netcdf split_file_2022121306-2022121310 {
dimensions:
	axis_nbounds = 2 ;
	lon = 1 ;
	lat = 1 ;
	nvertex = 2 ;
	levels = 39 ;
	time_counter = UNLIMITED ; // (5 currently)
variables:
	float lat(lat) ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:bounds = "bounds_lat" ;
	float lon(lon) ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:bounds = "bounds_lon" ;
	float bounds_lon(lat, lon, nvertex) ;
	float bounds_lat(lat, lon, nvertex) ;
	float levels(levels) ;
		levels:name = "levels" ;
		levels:units = "1" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 2022-12-13 01:00:00" ;
		time_instant:time_origin = "2022-12-13 01:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-12-13 01:00:00" ;
		time_counter:time_origin = "2022-12-13 01:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	float pressure(time_counter, levels, lat, lon) ;
		pressure:standard_name = "air_pressure" ;
		pressure:long_name = "Air Pressure" ;
		pressure:units = "Pa" ;
		pressure:online_operation = "instant" ;
		pressure:interval_operation = "1 h" ;
		pressure:interval_write = "1 h" ;
		pressure:cell_methods = "time: point" ;
		pressure:coordinates = "time_instant" ;
	float temperature(time_counter, levels, lat, lon) ;
		temperature:standard_name = "air_temperature" ;
		temperature:long_name = "Air Temperature" ;
		temperature:units = "K" ;
		temperature:online_operation = "instant" ;
		temperature:interval_operation = "1 h" ;
		temperature:interval_write = "1 h" ;
		temperature:cell_methods = "time: point" ;
		temperature:coordinates = "time_instant" ;

// global attributes:
		:name = "split_file" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "CF-1.6" ;
		:timeStamp = "2024-Jul-09 14:49:49 GMT" ;
		:uuid = "19159b97-0145-45c0-a68f-86e7ae916f0d" ;
data:

 lat = 51.5 ;

 lon = -4.5 ;

 bounds_lon =
  -6, -3 ;

 bounds_lat =
  50, 53 ;

 levels = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 171, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39 ;

 time_instant = 21600, 25200, 28800, 32400, 36000 ;

 time_instant_bounds =
  21600, 21600,
  25200, 25200,
  28800, 28800,
  32400, 32400,
  36000, 36000 ;

 time_counter = 21600, 25200, 28800, 32400, 36000 ;

 time_counter_bounds =
  21600, 21600,
  25200, 25200,
  28800, 28800,
  32400, 32400,
  36000, 36000 ;

 pressure =
  6099966,
  6099940,
  6099880,
  6099778,
  6099636,
  6099452,
  6099227,
  6098961,
  6098652,
  6098302,
  6097909,
  6097473,
  6096994,
  6096471,
  6095902,
  6095285,
  6094618,
  6093898,
  6093123,
  6092288,
  6091392,
  6090431,
  6089404,
  6088322,
  6087214,
  6086106,
  6085000,
  6083877,
  6082724,
  6081516,
  6080240,
  6078882,
  6077426,
  6075842,
  6074129,
  6072079,
  6069945,
  6065668,
  6063428,
  7099966,
  7099940,
  7099880,
  7099778,
  7099636,
  7099452,
  7099227,
  7098961,
  7098652,
  7098302,
  7097909,
  7097473,
  7096994,
  7096471,
  7095902,
  7095285,
  7094618,
  7093898,
  7093123,
  7092288,
  7091392,
  7090431,
  7089404,
  7088322,
  7087214,
  7086106,
  7085000,
  7083877,
  7082724,
  7081516,
  7080240,
  7078882,
  7077426,
  7075842,
  7074129,
  7072079,
  7069945,
  7065668,
  7063428,
  8099966,
  8099940,
  8099880,
  8099778,
  8099636,
  8099452,
  8099227,
  8098961,
  8098652,
  8098302,
  8097909,
  8097473,
  8096994,
  8096471,
  8095902,
  8095285,
  8094618,
  8093898,
  8093123,
  8092288,
  8091392,
  8090431,
  8089404,
  8088322,
  8087214,
  8086106,
  8085000,
  8083877,
  8082724,
  8081516,
  8080240,
  8078882,
  8077426,
  8075842,
  8074129,
  8072079,
  8069945,
  8065668,
  8063428,
  9099967,
  9099940,
  9099880,
  9099778,
  9099635,
  9099452,
  9099227,
  9098961,
  9098652,
  9098301,
  9097909,
  9097473,
  9096994,
  9096471,
  9095902,
  9095285,
  9094618,
  9093898,
  9093123,
  9092288,
  9091392,
  9090431,
  9089404,
  9088321,
  9087213,
  9086106,
  9084999,
  9083877,
  9082724,
  9081516,
  9080240,
  9078881,
  9077426,
  9075843,
  9074129,
  9072079,
  9069945,
  9065668,
  9063427,
  1.009997e+07,
  1.009994e+07,
  1.009988e+07,
  1.009978e+07,
  1.009964e+07,
  1.009945e+07,
  1.009923e+07,
  1.009896e+07,
  1.009865e+07,
  1.00983e+07,
  1.009791e+07,
  1.009747e+07,
  1.009699e+07,
  1.009647e+07,
  1.00959e+07,
  1.009528e+07,
  1.009462e+07,
  1.00939e+07,
  1.009312e+07,
  1.009229e+07,
  1.009139e+07,
  1.009043e+07,
  1.00894e+07,
  1.008832e+07,
  1.008721e+07,
  1.008611e+07,
  1.0085e+07,
  1.008388e+07,
  1.008272e+07,
  1.008152e+07,
  1.008024e+07,
  1.007888e+07,
  1.007743e+07,
  1.007584e+07,
  1.007413e+07,
  1.007208e+07,
  1.006994e+07,
  1.006567e+07,
  1.006343e+07 ;

 temperature =
  6000274,
  6000273,
  6000273,
  6000272,
  6000272,
  6000270,
  6000270,
  6000268,
  6000267,
  6000266,
  6000264,
  6000262,
  6000259,
  6000256,
  6000253,
  6000248,
  6000244,
  6000238,
  6000233,
  6000226,
  6000220,
  6000214,
  6000207,
  6000206,
  6000210,
  6000217,
  6000222,
  6000224,
  6000224,
  6000224,
  6000224,
  6000223,
  6000222,
  6000223,
  6000223,
  6000223,
  6000228,
  6000219,
  6000267,
  7000274,
  7000273,
  7000273,
  7000272,
  7000272,
  7000270,
  7000270,
  7000268,
  7000267,
  7000266,
  7000264,
  7000262,
  7000259,
  7000256,
  7000253,
  7000248,
  7000244,
  7000238,
  7000233,
  7000226,
  7000220,
  7000214,
  7000207,
  7000206,
  7000210,
  7000217,
  7000222,
  7000224,
  7000224,
  7000224,
  7000224,
  7000223,
  7000222,
  7000223,
  7000223,
  7000223,
  7000228,
  7000219,
  7000267,
  8000274,
  8000273,
  8000273,
  8000272,
  8000272,
  8000270,
  8000270,
  8000268,
  8000267,
  8000266,
  8000264,
  8000262,
  8000259,
  8000256,
  8000253,
  8000248,
  8000244,
  8000238,
  8000233,
  8000226,
  8000220,
  8000214,
  8000207,
  8000206,
  8000210,
  8000217,
  8000222,
  8000224,
  8000224,
  8000224,
  8000224,
  8000223,
  8000222,
  8000223,
  8000223,
  8000223,
  8000228,
  8000219,
  8000267,
  9000273,
  9000273,
  9000273,
  9000273,
  9000272,
  9000271,
  9000270,
  9000268,
  9000267,
  9000265,
  9000263,
  9000261,
  9000259,
  9000256,
  9000253,
  9000249,
  9000244,
  9000239,
  9000233,
  9000227,
  9000220,
  9000213,
  9000207,
  9000206,
  9000210,
  9000217,
  9000221,
  9000224,
  9000225,
  9000224,
  9000224,
  9000223,
  9000223,
  9000223,
  9000223,
  9000223,
  9000227,
  9000219,
  9000267,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000026e+07,
  1.000026e+07,
  1.000026e+07,
  1.000026e+07,
  1.000026e+07,
  1.000025e+07,
  1.000025e+07,
  1.000024e+07,
  1.000024e+07,
  1.000023e+07,
  1.000023e+07,
  1.000022e+07,
  1.000021e+07,
  1.000021e+07,
  1.000021e+07,
  1.000021e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000023e+07,
  1.000022e+07,
  1.000027e+07 ;
}
