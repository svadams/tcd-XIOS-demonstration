netcdf quant_bg_3_comp {
dimensions:
	x = 10 ;
	y = 10 ;
variables:
	float field(x, y) ;
		field:_QuantizeBitGroomNumberOfSignificantDigits = 3 ;
data:

 field =
  0, 0, 0, 0, 0, 0, -0, -5.738317e-42, -0, -5.738317e-42,
  0, 0.5878906, 0.9509277, 0.9511718, 0.5876465, 3.590685e-09, -0.5876465, 
    -0.9511718, -0.9509277, -0.5878906,
  0, 1.175781, 1.901855, 1.902344, 1.175293, 7.18137e-09, -1.175293, 
    -1.902344, -1.901855, -1.175781,
  0, 1.763672, 2.852539, 2.853515, 1.763184, 1.077205e-08, -1.763184, 
    -2.853515, -2.852539, -1.763672,
  0, 2.351562, 3.803711, 3.804687, 2.350586, 1.436274e-08, -2.350586, 
    -3.804687, -3.803711, -2.351562,
  0, 2.939453, 4.753906, 4.755859, 2.938477, 1.794979e-08, -2.938477, 
    -4.755859, -4.753906, -2.939453,
  0, 3.527344, 5.705078, 5.707031, 3.526367, 2.154411e-08, -3.526367, 
    -5.707031, -5.705078, -3.527344,
  0, 4.115234, 6.65625, 6.658203, 4.113281, 2.513116e-08, -4.113281, 
    -6.658203, -6.65625, -4.115234,
  0, 4.703125, 7.607422, 7.609375, 4.701172, 2.872548e-08, -4.701172, 
    -7.609375, -7.607422, -4.703125,
  0, 5.291015, 8.558594, 8.562499, 5.289062, 3.23198e-08, -5.289062, 
    -8.562499, -8.558594, -5.291015 ;
}
