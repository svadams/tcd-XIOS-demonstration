netcdf quant_gran_3_comp {
dimensions:
	x = 10 ;
	y = 10 ;
variables:
	float field(x, y) ;
		field:_QuantizeGranularBitRoundNumberOfSignificantDigits = 3 ;
data:

 field =
  0, 0, 0, 0, 0, 0, -0, -0, -0, -0,
  0, 0.5878906, 0.9511719, 0.9511719, 0.5878906, 3.587047e-09, -0.5878906, 
    -0.9511719, -0.9511719, -0.5878906,
  0, 1.171875, 1.898438, 1.898438, 1.171875, 7.18137e-09, -1.171875, 
    -1.898438, -1.898438, -1.171875,
  0, 1.765625, 2.851562, 2.851562, 1.765625, 1.076842e-08, -1.765625, 
    -2.851562, -2.851562, -1.765625,
  0, 2.351562, 3.804688, 3.804688, 2.351562, 1.437729e-08, -2.351562, 
    -3.804688, -3.804688, -2.351562,
  0, 2.9375, 4.757812, 4.757812, 2.9375, 1.792796e-08, -2.9375, -4.757812, 
    -4.757812, -2.9375,
  0, 3.523438, 5.703125, 5.703125, 3.523438, 2.153683e-08, -3.523438, 
    -5.703125, -5.703125, -3.523438,
  0, 4.117188, 6.65625, 6.65625, 4.117188, 2.514571e-08, -4.117188, -6.65625, 
    -6.65625, -4.117188,
  0, 4.703125, 7.609375, 7.609375, 4.703125, 2.869638e-08, -4.703125, 
    -7.609375, -7.609375, -4.703125,
  0, 5.289062, 8.5625, 8.5625, 5.289062, 3.230525e-08, -5.289062, -8.5625, 
    -8.5625, -5.289062 ;
}
