netcdf diag_file_2022121313-2022121316 {
dimensions:
	axis_nbounds = 2 ;
	lon = 1 ;
	lat = 1 ;
	nvertex = 2 ;
	levels = 39 ;
	time_counter = UNLIMITED ; // (1 currently)
variables:
	float lat(lat) ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:bounds = "bounds_lat" ;
	float lon(lon) ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:bounds = "bounds_lon" ;
	float bounds_lon(lat, lon, nvertex) ;
	float bounds_lat(lat, lon, nvertex) ;
	float levels(levels) ;
		levels:name = "levels" ;
		levels:units = "1" ;
	double time_centered(time_counter) ;
		time_centered:standard_name = "time" ;
		time_centered:long_name = "Time axis" ;
		time_centered:calendar = "gregorian" ;
		time_centered:units = "seconds since 2022-12-13 01:00:00" ;
		time_centered:time_origin = "2022-12-13 01:00:00" ;
		time_centered:bounds = "time_centered_bounds" ;
	double time_centered_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-12-13 01:00:00" ;
		time_counter:time_origin = "2022-12-13 01:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	float average_temperature(time_counter, levels, lat, lon) ;
		average_temperature:standard_name = "air_temperature" ;
		average_temperature:long_name = "Air Temperature" ;
		average_temperature:units = "K" ;
		average_temperature:online_operation = "average" ;
		average_temperature:interval_operation = "3 h" ;
		average_temperature:interval_write = "3 h" ;
		average_temperature:cell_methods = "time: mean" ;
		average_temperature:coordinates = "time_centered" ;

// global attributes:
		:name = "diag_file" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "CF-1.6" ;
		:timeStamp = "2025-Jun-17 07:58:53 GMT" ;
		:uuid = "5945a28c-5d4a-42df-a356-db9154d31057" ;
data:

 lat = 51.5 ;

 lon = -4.5 ;

 bounds_lon =
  -6, -3 ;

 bounds_lat =
  50, 53 ;

 levels = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 171, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39 ;

 time_centered = 48600 ;

 time_centered_bounds =
  43200, 54000 ;

 time_counter = 48600 ;

 time_counter_bounds =
  43200, 54000 ;

 average_temperature =
  287,
  282,
  277,
  272,
  267,
  262,
  257,
  252,
  247,
  242,
  237,
  232,
  227,
  222,
  217,
  212,
  207,
  202,
  197,
  192,
  187,
  182,
  177,
  172,
  167,
  162,
  157,
  152,
  147,
  142,
  137,
  132,
  127,
  122,
  117,
  112,
  107,
  102,
  97 ;
}
