netcdf split_file_2022121301-2022121305 {
dimensions:
	axis_nbounds = 2 ;
	lon = 1 ;
	lat = 1 ;
	nvertex = 2 ;
	levels = 39 ;
	time_counter = UNLIMITED ; // (5 currently)
variables:
	float lat(lat) ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:bounds = "bounds_lat" ;
	float lon(lon) ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:bounds = "bounds_lon" ;
	float bounds_lon(lat, lon, nvertex) ;
	float bounds_lat(lat, lon, nvertex) ;
	float levels(levels) ;
		levels:name = "levels" ;
		levels:units = "1" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 2022-12-13 01:00:00" ;
		time_instant:time_origin = "2022-12-13 01:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-12-13 01:00:00" ;
		time_counter:time_origin = "2022-12-13 01:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	float pressure(time_counter, levels, lat, lon) ;
		pressure:standard_name = "air_pressure" ;
		pressure:long_name = "Air Pressure" ;
		pressure:units = "Pa" ;
		pressure:online_operation = "instant" ;
		pressure:interval_operation = "1 h" ;
		pressure:interval_write = "1 h" ;
		pressure:cell_methods = "time: point" ;
		pressure:coordinates = "time_instant" ;
	float temperature(time_counter, levels, lat, lon) ;
		temperature:standard_name = "air_temperature" ;
		temperature:long_name = "Air Temperature" ;
		temperature:units = "K" ;
		temperature:online_operation = "instant" ;
		temperature:interval_operation = "1 h" ;
		temperature:interval_write = "1 h" ;
		temperature:cell_methods = "time: point" ;
		temperature:coordinates = "time_instant" ;

// global attributes:
		:name = "split_file" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "CF-1.6" ;
		:timeStamp = "2024-Jul-09 14:49:49 GMT" ;
		:uuid = "d2a21544-42d4-48e3-a960-137015dccc7d" ;
data:

 lat = 51.5 ;

 lon = -4.5 ;

 bounds_lon =
  -6, -3 ;

 bounds_lat =
  50, 53 ;

 levels = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 171, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39 ;

 time_instant = 3600, 7200, 10800, 14400, 18000 ;

 time_instant_bounds =
  3600, 3600,
  7200, 7200,
  10800, 10800,
  14400, 14400,
  18000, 18000 ;

 time_counter = 3600, 7200, 10800, 14400, 18000 ;

 time_counter_bounds =
  3600, 3600,
  7200, 7200,
  10800, 10800,
  14400, 14400,
  18000, 18000 ;

 pressure =
  1099966,
  1099940,
  1099880,
  1099778,
  1099635,
  1099452,
  1099227,
  1098961,
  1098652,
  1098302,
  1097909,
  1097473,
  1096994,
  1096471,
  1095902,
  1095285,
  1094618,
  1093898,
  1093123,
  1092288,
  1091392,
  1090431,
  1089404,
  1088321,
  1087213,
  1086106,
  1084999,
  1083877,
  1082724,
  1081516,
  1080240,
  1078881,
  1077426,
  1075842,
  1074129,
  1072079,
  1069945,
  1065668,
  1063427,
  2099966,
  2099940,
  2099880,
  2099778,
  2099635,
  2099452,
  2099227,
  2098961,
  2098652,
  2098302,
  2097909,
  2097473,
  2096994,
  2096471,
  2095902,
  2095285,
  2094618,
  2093898,
  2093123,
  2092288,
  2091392,
  2090431,
  2089404,
  2088321,
  2087213,
  2086106,
  2084999,
  2083877,
  2082724,
  2081516,
  2080240,
  2078881,
  2077426,
  2075842,
  2074129,
  2072079,
  2069945,
  2065668,
  2063427,
  3099966,
  3099940,
  3099880,
  3099778,
  3099635,
  3099452,
  3099227,
  3098961,
  3098652,
  3098302,
  3097909,
  3097473,
  3096994,
  3096471,
  3095902,
  3095285,
  3094618,
  3093898,
  3093123,
  3092288,
  3091392,
  3090431,
  3089404,
  3088322,
  3087214,
  3086106,
  3084999,
  3083877,
  3082724,
  3081516,
  3080240,
  3078881,
  3077426,
  3075842,
  3074129,
  3072079,
  3069945,
  3065668,
  3063427,
  4099966,
  4099940,
  4099880,
  4099778,
  4099635,
  4099452,
  4099227,
  4098961,
  4098652,
  4098302,
  4097909,
  4097473,
  4096994,
  4096471,
  4095902,
  4095285,
  4094618,
  4093898,
  4093123,
  4092288,
  4091392,
  4090431,
  4089404,
  4088322,
  4087214,
  4086106,
  4084999,
  4083877,
  4082724,
  4081516,
  4080240,
  4078881,
  4077426,
  4075842,
  4074129,
  4072079,
  4069945,
  4065668,
  4063427,
  5099966,
  5099940,
  5099880,
  5099778,
  5099636,
  5099452,
  5099227,
  5098961,
  5098652,
  5098302,
  5097909,
  5097473,
  5096994,
  5096471,
  5095902,
  5095285,
  5094618,
  5093898,
  5093123,
  5092288,
  5091392,
  5090431,
  5089404,
  5088322,
  5087214,
  5086106,
  5085000,
  5083877,
  5082724,
  5081516,
  5080240,
  5078882,
  5077426,
  5075842,
  5074129,
  5072079,
  5069945,
  5065668,
  5063428 ;

 temperature =
  1000273,
  1000273,
  1000273,
  1000272,
  1000272,
  1000271,
  1000270,
  1000268,
  1000267,
  1000265,
  1000263,
  1000262,
  1000259,
  1000256,
  1000253,
  1000249,
  1000244,
  1000239,
  1000233,
  1000227,
  1000220,
  1000214,
  1000207,
  1000206,
  1000210,
  1000217,
  1000221,
  1000224,
  1000225,
  1000224,
  1000224,
  1000223,
  1000223,
  1000223,
  1000223,
  1000223,
  1000227,
  1000219,
  1000267,
  2000273,
  2000273,
  2000273,
  2000272,
  2000272,
  2000271,
  2000270,
  2000268,
  2000267,
  2000265,
  2000263,
  2000262,
  2000259,
  2000256,
  2000253,
  2000249,
  2000244,
  2000239,
  2000233,
  2000227,
  2000220,
  2000214,
  2000207,
  2000206,
  2000210,
  2000217,
  2000222,
  2000224,
  2000225,
  2000224,
  2000224,
  2000223,
  2000223,
  2000223,
  2000223,
  2000223,
  2000227,
  2000219,
  2000267,
  3000274,
  3000273,
  3000273,
  3000272,
  3000272,
  3000271,
  3000270,
  3000268,
  3000267,
  3000265,
  3000264,
  3000262,
  3000259,
  3000256,
  3000253,
  3000249,
  3000244,
  3000238,
  3000233,
  3000227,
  3000220,
  3000214,
  3000207,
  3000206,
  3000210,
  3000217,
  3000222,
  3000224,
  3000225,
  3000224,
  3000224,
  3000223,
  3000223,
  3000223,
  3000223,
  3000223,
  3000227,
  3000219,
  3000267,
  4000274,
  4000273,
  4000273,
  4000272,
  4000272,
  4000271,
  4000270,
  4000268,
  4000267,
  4000265,
  4000264,
  4000262,
  4000259,
  4000256,
  4000253,
  4000249,
  4000244,
  4000238,
  4000233,
  4000227,
  4000220,
  4000214,
  4000207,
  4000206,
  4000210,
  4000217,
  4000222,
  4000224,
  4000225,
  4000224,
  4000224,
  4000223,
  4000223,
  4000223,
  4000223,
  4000223,
  4000227,
  4000219,
  4000267,
  5000274,
  5000273,
  5000273,
  5000272,
  5000272,
  5000270,
  5000270,
  5000268,
  5000267,
  5000266,
  5000264,
  5000262,
  5000259,
  5000256,
  5000253,
  5000248,
  5000244,
  5000238,
  5000233,
  5000226,
  5000220,
  5000214,
  5000207,
  5000206,
  5000210,
  5000217,
  5000222,
  5000224,
  5000224,
  5000224,
  5000224,
  5000223,
  5000222,
  5000223,
  5000223,
  5000223,
  5000228,
  5000219,
  5000267 ;
}
