netcdf reference_comp {
dimensions:
	x = 10 ;
	y = 10 ;
variables:
	float field(x, y) ;
data:

 field =
  0, 0, 0, 0, 0, 0, -0, -0, -0, -0,
  0, 0.5877852, 0.9510565, 0.9510565, 0.5877852, 3.589793e-09, -0.5877852, 
    -0.9510565, -0.9510565, -0.5877852,
  0, 1.17557, 1.902113, 1.902113, 1.17557, 7.179586e-09, -1.17557, -1.902113, 
    -1.902113, -1.17557,
  0, 1.763356, 2.853169, 2.853169, 1.763356, 1.076938e-08, -1.763356, 
    -2.853169, -2.853169, -1.763356,
  0, 2.351141, 3.804226, 3.804226, 2.351141, 1.435917e-08, -2.351141, 
    -3.804226, -3.804226, -2.351141,
  0, 2.938926, 4.755282, 4.755282, 2.938926, 1.794896e-08, -2.938926, 
    -4.755282, -4.755282, -2.938926,
  0, 3.526711, 5.706339, 5.706339, 3.526711, 2.153876e-08, -3.526711, 
    -5.706339, -5.706339, -3.526711,
  0, 4.114497, 6.657396, 6.657396, 4.114497, 2.512855e-08, -4.114497, 
    -6.657396, -6.657396, -4.114497,
  0, 4.702282, 7.608452, 7.608452, 4.702282, 2.871835e-08, -4.702282, 
    -7.608452, -7.608452, -4.702282,
  0, 5.290067, 8.559508, 8.559508, 5.290067, 3.230814e-08, -5.290067, 
    -8.559508, -8.559508, -5.290067 ;
}
