netcdf mixed_frequency {
dimensions:
	axis_nbounds = 2 ;
	lon = 1 ;
	lat = 1 ;
	nvertex = 2 ;
	levels = 39 ;
	time_counter = UNLIMITED ; // (20 currently)
variables:
	float lat(lat) ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:bounds = "bounds_lat" ;
	float lon(lon) ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:bounds = "bounds_lon" ;
	float bounds_lon(lat, lon, nvertex) ;
	float bounds_lat(lat, lon, nvertex) ;
	float levels(levels) ;
		levels:name = "levels" ;
		levels:units = "1" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 2022-12-13 01:00:00" ;
		time_instant:time_origin = "2022-12-13 01:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-12-13 01:00:00" ;
		time_counter:time_origin = "2022-12-13 01:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	float pressure(time_counter, levels, lat, lon) ;
		pressure:standard_name = "air_pressure" ;
		pressure:long_name = "Air Pressure" ;
		pressure:units = "Pa" ;
		pressure:online_operation = "instant" ;
		pressure:interval_operation = "1 h" ;
		pressure:interval_write = "1 h" ;
		pressure:cell_methods = "time: point" ;
		pressure:coordinates = "time_instant" ;
	float temperature(time_counter, levels, lat, lon) ;
		temperature:standard_name = "air_temperature" ;
		temperature:long_name = "Air Temperature" ;
		temperature:units = "K" ;
		temperature:online_operation = "instant" ;
		temperature:interval_operation = "1 h" ;
		temperature:interval_write = "1 h" ;
		temperature:cell_methods = "time: point" ;
		temperature:coordinates = "time_instant" ;

// global attributes:
		:name = "mixed_frequency" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "CF-1.6" ;
		:timeStamp = "2024-Jul-09 10:21:42 GMT" ;
		:uuid = "6f3f15c1-40e6-481b-9d82-af0d1524fe5e" ;
data:

 lat = 51.5 ;

 lon = -4.5 ;

 bounds_lon =
  -6, -3 ;

 bounds_lat =
  50, 53 ;

 levels = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 171, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39 ;

 time_instant = 3600, 7200, 10800, 14400, 18000, 21600, 25200, 28800, 32400, 
    36000, 39600, 43200, 46800, 50400, 54000, 57600, 61200, 64800, 68400, 
    72000 ;

 time_instant_bounds =
  3600, 3600,
  7200, 7200,
  10800, 10800,
  14400, 14400,
  18000, 18000,
  21600, 21600,
  25200, 25200,
  28800, 28800,
  32400, 32400,
  36000, 36000,
  39600, 39600,
  43200, 43200,
  46800, 46800,
  50400, 50400,
  54000, 54000,
  57600, 57600,
  61200, 61200,
  64800, 64800,
  68400, 68400,
  72000, 72000 ;

 time_counter = 3600, 7200, 10800, 14400, 18000, 21600, 25200, 28800, 32400, 
    36000, 39600, 43200, 46800, 50400, 54000, 57600, 61200, 64800, 68400, 
    72000 ;

 time_counter_bounds =
  3600, 3600,
  7200, 7200,
  10800, 10800,
  14400, 14400,
  18000, 18000,
  21600, 21600,
  25200, 25200,
  28800, 28800,
  32400, 32400,
  36000, 36000,
  39600, 39600,
  43200, 43200,
  46800, 46800,
  50400, 50400,
  54000, 54000,
  57600, 57600,
  61200, 61200,
  64800, 64800,
  68400, 68400,
  72000, 72000 ;

 pressure =
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  3099966,
  3099940,
  3099880,
  3099778,
  3099635,
  3099452,
  3099227,
  3098961,
  3098652,
  3098302,
  3097909,
  3097473,
  3096994,
  3096471,
  3095902,
  3095285,
  3094618,
  3093898,
  3093123,
  3092288,
  3091392,
  3090431,
  3089404,
  3088322,
  3087214,
  3086106,
  3084999,
  3083877,
  3082724,
  3081516,
  3080240,
  3078881,
  3077426,
  3075842,
  3074129,
  3072079,
  3069945,
  3065668,
  3063427,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  6099966,
  6099940,
  6099880,
  6099778,
  6099636,
  6099452,
  6099227,
  6098961,
  6098652,
  6098302,
  6097909,
  6097473,
  6096994,
  6096471,
  6095902,
  6095285,
  6094618,
  6093898,
  6093123,
  6092288,
  6091392,
  6090431,
  6089404,
  6088322,
  6087214,
  6086106,
  6085000,
  6083877,
  6082724,
  6081516,
  6080240,
  6078882,
  6077426,
  6075842,
  6074129,
  6072079,
  6069945,
  6065668,
  6063428,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  9099967,
  9099940,
  9099880,
  9099778,
  9099635,
  9099452,
  9099227,
  9098961,
  9098652,
  9098301,
  9097909,
  9097473,
  9096994,
  9096471,
  9095902,
  9095285,
  9094618,
  9093898,
  9093123,
  9092288,
  9091392,
  9090431,
  9089404,
  9088321,
  9087213,
  9086106,
  9084999,
  9083877,
  9082724,
  9081516,
  9080240,
  9078881,
  9077426,
  9075843,
  9074129,
  9072079,
  9069945,
  9065668,
  9063427,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.209997e+07,
  1.209994e+07,
  1.209988e+07,
  1.209978e+07,
  1.209964e+07,
  1.209945e+07,
  1.209923e+07,
  1.209896e+07,
  1.209865e+07,
  1.20983e+07,
  1.209791e+07,
  1.209747e+07,
  1.209699e+07,
  1.209647e+07,
  1.20959e+07,
  1.209528e+07,
  1.209462e+07,
  1.20939e+07,
  1.209312e+07,
  1.209229e+07,
  1.209139e+07,
  1.209043e+07,
  1.20894e+07,
  1.208832e+07,
  1.208721e+07,
  1.208611e+07,
  1.2085e+07,
  1.208388e+07,
  1.208272e+07,
  1.208152e+07,
  1.208024e+07,
  1.207888e+07,
  1.207743e+07,
  1.207584e+07,
  1.207413e+07,
  1.207208e+07,
  1.206994e+07,
  1.206567e+07,
  1.206343e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.509997e+07,
  1.509994e+07,
  1.509988e+07,
  1.509978e+07,
  1.509964e+07,
  1.509945e+07,
  1.509923e+07,
  1.509896e+07,
  1.509865e+07,
  1.50983e+07,
  1.509791e+07,
  1.509747e+07,
  1.509699e+07,
  1.509647e+07,
  1.50959e+07,
  1.509528e+07,
  1.509462e+07,
  1.50939e+07,
  1.509312e+07,
  1.509229e+07,
  1.509139e+07,
  1.509043e+07,
  1.50894e+07,
  1.508832e+07,
  1.508721e+07,
  1.508611e+07,
  1.5085e+07,
  1.508388e+07,
  1.508272e+07,
  1.508152e+07,
  1.508024e+07,
  1.507888e+07,
  1.507743e+07,
  1.507584e+07,
  1.507413e+07,
  1.507208e+07,
  1.506994e+07,
  1.506567e+07,
  1.506343e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.809997e+07,
  1.809994e+07,
  1.809988e+07,
  1.809978e+07,
  1.809964e+07,
  1.809945e+07,
  1.809923e+07,
  1.809896e+07,
  1.809865e+07,
  1.80983e+07,
  1.809791e+07,
  1.809747e+07,
  1.809699e+07,
  1.809647e+07,
  1.80959e+07,
  1.809528e+07,
  1.809462e+07,
  1.80939e+07,
  1.809312e+07,
  1.809229e+07,
  1.809139e+07,
  1.809043e+07,
  1.80894e+07,
  1.808832e+07,
  1.808721e+07,
  1.808611e+07,
  1.8085e+07,
  1.808388e+07,
  1.808272e+07,
  1.808152e+07,
  1.808024e+07,
  1.807888e+07,
  1.807743e+07,
  1.807584e+07,
  1.807413e+07,
  1.807208e+07,
  1.806995e+07,
  1.806567e+07,
  1.806343e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _ ;

 temperature =
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  2000273,
  2000273,
  2000273,
  2000272,
  2000272,
  2000271,
  2000270,
  2000268,
  2000267,
  2000265,
  2000263,
  2000262,
  2000259,
  2000256,
  2000253,
  2000249,
  2000244,
  2000239,
  2000233,
  2000227,
  2000220,
  2000214,
  2000207,
  2000206,
  2000210,
  2000217,
  2000222,
  2000224,
  2000225,
  2000224,
  2000224,
  2000223,
  2000223,
  2000223,
  2000223,
  2000223,
  2000227,
  2000219,
  2000267,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  4000274,
  4000273,
  4000273,
  4000272,
  4000272,
  4000271,
  4000270,
  4000268,
  4000267,
  4000265,
  4000264,
  4000262,
  4000259,
  4000256,
  4000253,
  4000249,
  4000244,
  4000238,
  4000233,
  4000227,
  4000220,
  4000214,
  4000207,
  4000206,
  4000210,
  4000217,
  4000222,
  4000224,
  4000225,
  4000224,
  4000224,
  4000223,
  4000223,
  4000223,
  4000223,
  4000223,
  4000227,
  4000219,
  4000267,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  6000274,
  6000273,
  6000273,
  6000272,
  6000272,
  6000270,
  6000270,
  6000268,
  6000267,
  6000266,
  6000264,
  6000262,
  6000259,
  6000256,
  6000253,
  6000248,
  6000244,
  6000238,
  6000233,
  6000226,
  6000220,
  6000214,
  6000207,
  6000206,
  6000210,
  6000217,
  6000222,
  6000224,
  6000224,
  6000224,
  6000224,
  6000223,
  6000222,
  6000223,
  6000223,
  6000223,
  6000228,
  6000219,
  6000267,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  8000274,
  8000273,
  8000273,
  8000272,
  8000272,
  8000270,
  8000270,
  8000268,
  8000267,
  8000266,
  8000264,
  8000262,
  8000259,
  8000256,
  8000253,
  8000248,
  8000244,
  8000238,
  8000233,
  8000226,
  8000220,
  8000214,
  8000207,
  8000206,
  8000210,
  8000217,
  8000222,
  8000224,
  8000224,
  8000224,
  8000224,
  8000223,
  8000222,
  8000223,
  8000223,
  8000223,
  8000228,
  8000219,
  8000267,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000027e+07,
  1.000026e+07,
  1.000026e+07,
  1.000026e+07,
  1.000026e+07,
  1.000026e+07,
  1.000025e+07,
  1.000025e+07,
  1.000024e+07,
  1.000024e+07,
  1.000023e+07,
  1.000023e+07,
  1.000022e+07,
  1.000021e+07,
  1.000021e+07,
  1.000021e+07,
  1.000021e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000022e+07,
  1.000023e+07,
  1.000022e+07,
  1.000027e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200026e+07,
  1.200026e+07,
  1.200026e+07,
  1.200026e+07,
  1.200026e+07,
  1.200025e+07,
  1.200025e+07,
  1.200024e+07,
  1.200024e+07,
  1.200023e+07,
  1.200023e+07,
  1.200022e+07,
  1.200021e+07,
  1.200021e+07,
  1.200021e+07,
  1.200021e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200023e+07,
  1.200022e+07,
  1.200027e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400026e+07,
  1.400026e+07,
  1.400026e+07,
  1.400026e+07,
  1.400026e+07,
  1.400025e+07,
  1.400025e+07,
  1.400024e+07,
  1.400024e+07,
  1.400023e+07,
  1.400023e+07,
  1.400022e+07,
  1.400021e+07,
  1.400021e+07,
  1.400021e+07,
  1.400021e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400023e+07,
  1.400022e+07,
  1.400027e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600026e+07,
  1.600026e+07,
  1.600026e+07,
  1.600026e+07,
  1.600026e+07,
  1.600025e+07,
  1.600025e+07,
  1.600024e+07,
  1.600024e+07,
  1.600023e+07,
  1.600023e+07,
  1.600022e+07,
  1.600021e+07,
  1.600021e+07,
  1.600021e+07,
  1.600021e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600023e+07,
  1.600022e+07,
  1.600027e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800026e+07,
  1.800026e+07,
  1.800026e+07,
  1.800026e+07,
  1.800025e+07,
  1.800025e+07,
  1.800024e+07,
  1.800024e+07,
  1.800023e+07,
  1.800023e+07,
  1.800022e+07,
  1.800021e+07,
  1.800021e+07,
  1.800021e+07,
  1.800021e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800023e+07,
  1.800022e+07,
  1.800027e+07,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  _,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000026e+07,
  2.000026e+07,
  2.000026e+07,
  2.000026e+07,
  2.000025e+07,
  2.000025e+07,
  2.000024e+07,
  2.000024e+07,
  2.000023e+07,
  2.000023e+07,
  2.000022e+07,
  2.000021e+07,
  2.000021e+07,
  2.000021e+07,
  2.000021e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000023e+07,
  2.000022e+07,
  2.000027e+07 ;
}
