netcdf quant_br_10b_comp {
dimensions:
	x = 10 ;
	y = 10 ;
variables:
	float field(x, y) ;
		field:_QuantizeBitRoundNumberOfSignificantBits = 10 ;
data:

 field =
  0, 0, 0, 0, 0, 0, -0, -0, -0, -0,
  0, 0.5878906, 0.9511719, 0.9511719, 0.5878906, 3.590685e-09, -0.5878906, 
    -0.9511719, -0.9511719, -0.5878906,
  0, 1.175781, 1.902344, 1.902344, 1.175781, 7.18137e-09, -1.175781, 
    -1.902344, -1.902344, -1.175781,
  0, 1.763672, 2.853516, 2.853516, 1.763672, 1.076842e-08, -1.763672, 
    -2.853516, -2.853516, -1.763672,
  0, 2.351562, 3.804688, 3.804688, 2.351562, 1.436274e-08, -2.351562, 
    -3.804688, -3.804688, -2.351562,
  0, 2.939453, 4.753906, 4.753906, 2.939453, 1.794251e-08, -2.939453, 
    -4.753906, -4.753906, -2.939453,
  0, 3.527344, 5.707031, 5.707031, 3.527344, 2.153683e-08, -3.527344, 
    -5.707031, -5.707031, -3.527344,
  0, 4.113281, 6.65625, 6.65625, 4.113281, 2.513116e-08, -4.113281, -6.65625, 
    -6.65625, -4.113281,
  0, 4.703125, 7.609375, 7.609375, 4.703125, 2.872548e-08, -4.703125, 
    -7.609375, -7.609375, -4.703125,
  0, 5.289062, 8.5625, 8.5625, 5.289062, 3.230525e-08, -5.289062, -8.5625, 
    -8.5625, -5.289062 ;
}
