netcdf split_file_2022121311-2022121315 {
dimensions:
	axis_nbounds = 2 ;
	lon = 1 ;
	lat = 1 ;
	nvertex = 2 ;
	levels = 39 ;
	time_counter = UNLIMITED ; // (5 currently)
variables:
	float lat(lat) ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:bounds = "bounds_lat" ;
	float lon(lon) ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:bounds = "bounds_lon" ;
	float bounds_lon(lat, lon, nvertex) ;
	float bounds_lat(lat, lon, nvertex) ;
	float levels(levels) ;
		levels:name = "levels" ;
		levels:units = "1" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 2022-12-13 01:00:00" ;
		time_instant:time_origin = "2022-12-13 01:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-12-13 01:00:00" ;
		time_counter:time_origin = "2022-12-13 01:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	float pressure(time_counter, levels, lat, lon) ;
		pressure:standard_name = "air_pressure" ;
		pressure:long_name = "Air Pressure" ;
		pressure:units = "Pa" ;
		pressure:online_operation = "instant" ;
		pressure:interval_operation = "1 h" ;
		pressure:interval_write = "1 h" ;
		pressure:cell_methods = "time: point" ;
		pressure:coordinates = "time_instant" ;
	float temperature(time_counter, levels, lat, lon) ;
		temperature:standard_name = "air_temperature" ;
		temperature:long_name = "Air Temperature" ;
		temperature:units = "K" ;
		temperature:online_operation = "instant" ;
		temperature:interval_operation = "1 h" ;
		temperature:interval_write = "1 h" ;
		temperature:cell_methods = "time: point" ;
		temperature:coordinates = "time_instant" ;

// global attributes:
		:name = "split_file" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "CF-1.6" ;
		:timeStamp = "2024-Jul-09 14:49:49 GMT" ;
		:uuid = "895bd342-97e4-4a74-8396-18394e7c07ab" ;
data:

 lat = 51.5 ;

 lon = -4.5 ;

 bounds_lon =
  -6, -3 ;

 bounds_lat =
  50, 53 ;

 levels = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 171, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39 ;

 time_instant = 39600, 43200, 46800, 50400, 54000 ;

 time_instant_bounds =
  39600, 39600,
  43200, 43200,
  46800, 46800,
  50400, 50400,
  54000, 54000 ;

 time_counter = 39600, 43200, 46800, 50400, 54000 ;

 time_counter_bounds =
  39600, 39600,
  43200, 43200,
  46800, 46800,
  50400, 50400,
  54000, 54000 ;

 pressure =
  1.109997e+07,
  1.109994e+07,
  1.109988e+07,
  1.109978e+07,
  1.109964e+07,
  1.109945e+07,
  1.109923e+07,
  1.109896e+07,
  1.109865e+07,
  1.10983e+07,
  1.109791e+07,
  1.109747e+07,
  1.109699e+07,
  1.109647e+07,
  1.10959e+07,
  1.109528e+07,
  1.109462e+07,
  1.10939e+07,
  1.109312e+07,
  1.109229e+07,
  1.109139e+07,
  1.109043e+07,
  1.10894e+07,
  1.108832e+07,
  1.108721e+07,
  1.108611e+07,
  1.1085e+07,
  1.108388e+07,
  1.108272e+07,
  1.108152e+07,
  1.108024e+07,
  1.107888e+07,
  1.107743e+07,
  1.107584e+07,
  1.107413e+07,
  1.107208e+07,
  1.106994e+07,
  1.106567e+07,
  1.106343e+07,
  1.209997e+07,
  1.209994e+07,
  1.209988e+07,
  1.209978e+07,
  1.209964e+07,
  1.209945e+07,
  1.209923e+07,
  1.209896e+07,
  1.209865e+07,
  1.20983e+07,
  1.209791e+07,
  1.209747e+07,
  1.209699e+07,
  1.209647e+07,
  1.20959e+07,
  1.209528e+07,
  1.209462e+07,
  1.20939e+07,
  1.209312e+07,
  1.209229e+07,
  1.209139e+07,
  1.209043e+07,
  1.20894e+07,
  1.208832e+07,
  1.208721e+07,
  1.208611e+07,
  1.2085e+07,
  1.208388e+07,
  1.208272e+07,
  1.208152e+07,
  1.208024e+07,
  1.207888e+07,
  1.207743e+07,
  1.207584e+07,
  1.207413e+07,
  1.207208e+07,
  1.206994e+07,
  1.206567e+07,
  1.206343e+07,
  1.309997e+07,
  1.309994e+07,
  1.309988e+07,
  1.309978e+07,
  1.309964e+07,
  1.309945e+07,
  1.309923e+07,
  1.309896e+07,
  1.309865e+07,
  1.30983e+07,
  1.309791e+07,
  1.309747e+07,
  1.309699e+07,
  1.309647e+07,
  1.30959e+07,
  1.309528e+07,
  1.309462e+07,
  1.30939e+07,
  1.309312e+07,
  1.309229e+07,
  1.309139e+07,
  1.309043e+07,
  1.30894e+07,
  1.308832e+07,
  1.308721e+07,
  1.308611e+07,
  1.3085e+07,
  1.308388e+07,
  1.308272e+07,
  1.308152e+07,
  1.308024e+07,
  1.307888e+07,
  1.307743e+07,
  1.307584e+07,
  1.307413e+07,
  1.307208e+07,
  1.306994e+07,
  1.306567e+07,
  1.306343e+07,
  1.409997e+07,
  1.409994e+07,
  1.409988e+07,
  1.409978e+07,
  1.409964e+07,
  1.409945e+07,
  1.409923e+07,
  1.409896e+07,
  1.409865e+07,
  1.40983e+07,
  1.409791e+07,
  1.409747e+07,
  1.409699e+07,
  1.409647e+07,
  1.40959e+07,
  1.409528e+07,
  1.409462e+07,
  1.40939e+07,
  1.409312e+07,
  1.409229e+07,
  1.409139e+07,
  1.409043e+07,
  1.40894e+07,
  1.408832e+07,
  1.408721e+07,
  1.408611e+07,
  1.4085e+07,
  1.408388e+07,
  1.408272e+07,
  1.408152e+07,
  1.408024e+07,
  1.407888e+07,
  1.407743e+07,
  1.407584e+07,
  1.407413e+07,
  1.407208e+07,
  1.406994e+07,
  1.406567e+07,
  1.406343e+07,
  1.509997e+07,
  1.509994e+07,
  1.509988e+07,
  1.509978e+07,
  1.509964e+07,
  1.509945e+07,
  1.509923e+07,
  1.509896e+07,
  1.509865e+07,
  1.50983e+07,
  1.509791e+07,
  1.509747e+07,
  1.509699e+07,
  1.509647e+07,
  1.50959e+07,
  1.509528e+07,
  1.509462e+07,
  1.50939e+07,
  1.509312e+07,
  1.509229e+07,
  1.509139e+07,
  1.509043e+07,
  1.50894e+07,
  1.508832e+07,
  1.508721e+07,
  1.508611e+07,
  1.5085e+07,
  1.508388e+07,
  1.508272e+07,
  1.508152e+07,
  1.508024e+07,
  1.507888e+07,
  1.507743e+07,
  1.507584e+07,
  1.507413e+07,
  1.507208e+07,
  1.506994e+07,
  1.506567e+07,
  1.506343e+07 ;

 temperature =
  1.100027e+07,
  1.100027e+07,
  1.100027e+07,
  1.100027e+07,
  1.100027e+07,
  1.100027e+07,
  1.100027e+07,
  1.100027e+07,
  1.100027e+07,
  1.100026e+07,
  1.100026e+07,
  1.100026e+07,
  1.100026e+07,
  1.100026e+07,
  1.100025e+07,
  1.100025e+07,
  1.100024e+07,
  1.100024e+07,
  1.100023e+07,
  1.100023e+07,
  1.100022e+07,
  1.100021e+07,
  1.100021e+07,
  1.100021e+07,
  1.100021e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100022e+07,
  1.100023e+07,
  1.100022e+07,
  1.100027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200027e+07,
  1.200026e+07,
  1.200026e+07,
  1.200026e+07,
  1.200026e+07,
  1.200026e+07,
  1.200025e+07,
  1.200025e+07,
  1.200024e+07,
  1.200024e+07,
  1.200023e+07,
  1.200023e+07,
  1.200022e+07,
  1.200021e+07,
  1.200021e+07,
  1.200021e+07,
  1.200021e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200022e+07,
  1.200023e+07,
  1.200022e+07,
  1.200027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300027e+07,
  1.300026e+07,
  1.300026e+07,
  1.300026e+07,
  1.300026e+07,
  1.300026e+07,
  1.300025e+07,
  1.300025e+07,
  1.300024e+07,
  1.300024e+07,
  1.300023e+07,
  1.300023e+07,
  1.300022e+07,
  1.300021e+07,
  1.300021e+07,
  1.300021e+07,
  1.300021e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300022e+07,
  1.300023e+07,
  1.300022e+07,
  1.300027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400027e+07,
  1.400026e+07,
  1.400026e+07,
  1.400026e+07,
  1.400026e+07,
  1.400026e+07,
  1.400025e+07,
  1.400025e+07,
  1.400024e+07,
  1.400024e+07,
  1.400023e+07,
  1.400023e+07,
  1.400022e+07,
  1.400021e+07,
  1.400021e+07,
  1.400021e+07,
  1.400021e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400022e+07,
  1.400023e+07,
  1.400022e+07,
  1.400027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500027e+07,
  1.500026e+07,
  1.500026e+07,
  1.500026e+07,
  1.500026e+07,
  1.500026e+07,
  1.500025e+07,
  1.500025e+07,
  1.500024e+07,
  1.500024e+07,
  1.500023e+07,
  1.500023e+07,
  1.500022e+07,
  1.500021e+07,
  1.500021e+07,
  1.500021e+07,
  1.500021e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500022e+07,
  1.500023e+07,
  1.500022e+07,
  1.500027e+07 ;
}
