netcdf domain_input {
dimensions:
        x = 5 ;
        y = 5 ;
        x_resample = 2 ;
        y_resample = 2 ;
variables:
        float x(x) ;
                x:long_name = "original x coordinate" ;
                x:units = "1";
        float y(y) ;
                y:long_name = "original y coordinate" ;
                y:units = "1";
        float x_resample(x_resample) ;
                x_resample:long_name = "resampled x coordinate" ;
                x_resample:units = "1";
        float y_resample(y_resample) ;
                y_resample:long_name = "resampled y coordinate" ;
                y_resample:units = "1";
        double original_data(y,x) ;
                original_data:long_name = "input data values" ;
                original_data:units = "1";
        double resample_data(y_resample,x_resample) ;
                resample_data:long_name = "expected resampled data values" ;
                resample_data:units = "1";

// global attributes:
                :title = "Input data for XIOS Domain resampling; data is a square function of the x & y coordinates; x^2+y^2." ;

data:

 x = 0, 2, 4, 6, 8 ;

 y = 0, 2, 4, 6, 8 ;

 x_resample = 3, 5 ;

 y_resample = 3, 5 ;

 original_data =  0,  4, 16, 36, 64,
                  4,  8, 20, 40, 68,
                 16, 20, 32, 52, 80,
                 36, 40, 52, 72, 100,
                 64, 68, 80, 100, 128 ;

 resample_data = 18, 34,
                 34, 50 ;

}
