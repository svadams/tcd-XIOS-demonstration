netcdf input_2 {
dimensions:
	axis_nbounds = 2 ;
	lon = 2 ;
	lat = 2 ;
	model_axis = 1 ;
	time_counter = UNLIMITED ; // (1 currently)
variables:
	float model_axis(model_axis) ;
		model_axis:name = "model_axis" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "360_day" ;
		time_instant:units = "seconds since 2012-02-29 15:00:00" ;
		time_instant:time_origin = "2012-02-29 15:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "360_day" ;
		time_counter:units = "seconds since 2012-02-29 15:00:00" ;
		time_counter:time_origin = "2012-02-29 15:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	float field_B(time_counter, model_axis, lat, lon) ;
		field_B:online_operation = "instant" ;
		field_B:interval_operation = "1 h" ;
		field_B:interval_write = "1 h" ;
		field_B:cell_methods = "time: point" ;
		field_B:coordinates = "time_instant" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.10.0" ;
		:name = "input_2" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "CF-1.6" ;
		:timeStamp = "2024-Apr-23 16:06:49 GMT" ;
		:uuid = "7ed89cad-d456-41f0-8e3b-b4fb817d68fd" ;
data:

 model_axis = 1 ;

 time_instant = 176400 ;

 time_instant_bounds =
  176400, 176400 ;

 time_counter = 176400 ;

 time_counter_bounds =
  176400, 176400 ;

 field_B =
  1, 1,
  1, 1 ;
}
