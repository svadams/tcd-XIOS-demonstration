netcdf mesh_C12 {
dimensions:
	ndynamics_node = 866 ;
	ndynamics_edge = 1728 ;
	ndynamics_face = 864 ;
	One = 1 ;
	Two = 2 ;
	Four = 4 ;
variables:
	int dynamics ;
		dynamics:cf_role = "mesh_topology" ;
		dynamics:geometry = "spherical" ;
		dynamics:topology = "periodic" ;
		dynamics:coord_sys = "ll" ;
		dynamics:max_stencil_depth = 0 ;
		dynamics:periodic_x = "F" ;
		dynamics:periodic_y = "F" ;
		dynamics:constructor_inputs = "edge_cells=12;smooth_passes=0" ;
		dynamics:n_mesh_maps = 0 ;
		dynamics:long_name = "Topology data of 2D unstructured mesh" ;
		dynamics:topology_dimension = 2 ;
		dynamics:node_coordinates = "dynamics_node_x dynamics_node_y" ;
		dynamics:face_coordinates = "dynamics_face_x dynamics_face_y" ;
		dynamics:face_node_connectivity = "dynamics_face_nodes" ;
		dynamics:edge_node_connectivity = "dynamics_edge_nodes" ;
		dynamics:face_edge_connectivity = "dynamics_face_edges" ;
		dynamics:face_face_connectivity = "dynamics_face_links" ;
		dynamics:north_pole = 0., 90. ;
		dynamics:null_island = 0., 0. ;
	int dynamics_face_nodes(ndynamics_face, Four) ;
		dynamics_face_nodes:cf_role = "face_node_connectivity" ;
		dynamics_face_nodes:long_name = "Maps every quadrilateral face to its four corner nodes." ;
		dynamics_face_nodes:start_index = 1 ;
	int dynamics_edge_nodes(ndynamics_edge, Two) ;
		dynamics_edge_nodes:cf_role = "edge_node_connectivity" ;
		dynamics_edge_nodes:long_name = "Maps every edge to the two nodes that it connects." ;
		dynamics_edge_nodes:start_index = 1 ;
	int dynamics_face_edges(ndynamics_face, Four) ;
		dynamics_face_edges:cf_role = "face_edge_connectivity" ;
		dynamics_face_edges:long_name = "Maps every quadrilateral face to its four edges." ;
		dynamics_face_edges:start_index = 1 ;
	int dynamics_face_links(ndynamics_face, Four) ;
		dynamics_face_links:cf_role = "face_face_connectivity" ;
		dynamics_face_links:long_name = "Indicates which other faces neighbour each face." ;
		dynamics_face_links:start_index = 1 ;
		dynamics_face_links:flag_values = -1 ;
		dynamics_face_links:flag_meanings = "out_of_mesh" ;
	double dynamics_node_x(ndynamics_node) ;
		dynamics_node_x:standard_name = "longitude" ;
		dynamics_node_x:long_name = "longitude of 2D mesh nodes." ;
		dynamics_node_x:units = "degrees_east" ;
	double dynamics_node_y(ndynamics_node) ;
		dynamics_node_y:standard_name = "latitude" ;
		dynamics_node_y:long_name = "latitude of 2D mesh nodes." ;
		dynamics_node_y:units = "degrees_north" ;
	double dynamics_face_x(ndynamics_face) ;
		dynamics_face_x:standard_name = "longitude" ;
		dynamics_face_x:long_name = "longitude of 2D face centres" ;
		dynamics_face_x:units = "degrees_east" ;
	double dynamics_face_y(ndynamics_face) ;
		dynamics_face_y:standard_name = "latitude" ;
		dynamics_face_y:long_name = "latitude of 2D face centres" ;
		dynamics_face_y:units = "degrees_north" ;
data:

 dynamics = _ ;

 dynamics_face_nodes =
  13, 14, 2, 1,
  14, 15, 3, 2,
  15, 16, 4, 3,
  16, 17, 5, 4,
  17, 18, 6, 5,
  18, 19, 7, 6,
  19, 20, 8, 7,
  20, 21, 9, 8,
  21, 22, 10, 9,
  22, 23, 11, 10,
  23, 24, 12, 11,
  24, 157, 145, 12,
  25, 26, 14, 13,
  26, 27, 15, 14,
  27, 28, 16, 15,
  28, 29, 17, 16,
  29, 30, 18, 17,
  30, 31, 19, 18,
  31, 32, 20, 19,
  32, 33, 21, 20,
  33, 34, 22, 21,
  34, 35, 23, 22,
  35, 36, 24, 23,
  36, 169, 157, 24,
  37, 38, 26, 25,
  38, 39, 27, 26,
  39, 40, 28, 27,
  40, 41, 29, 28,
  41, 42, 30, 29,
  42, 43, 31, 30,
  43, 44, 32, 31,
  44, 45, 33, 32,
  45, 46, 34, 33,
  46, 47, 35, 34,
  47, 48, 36, 35,
  48, 181, 169, 36,
  49, 50, 38, 37,
  50, 51, 39, 38,
  51, 52, 40, 39,
  52, 53, 41, 40,
  53, 54, 42, 41,
  54, 55, 43, 42,
  55, 56, 44, 43,
  56, 57, 45, 44,
  57, 58, 46, 45,
  58, 59, 47, 46,
  59, 60, 48, 47,
  60, 193, 181, 48,
  61, 62, 50, 49,
  62, 63, 51, 50,
  63, 64, 52, 51,
  64, 65, 53, 52,
  65, 66, 54, 53,
  66, 67, 55, 54,
  67, 68, 56, 55,
  68, 69, 57, 56,
  69, 70, 58, 57,
  70, 71, 59, 58,
  71, 72, 60, 59,
  72, 205, 193, 60,
  73, 74, 62, 61,
  74, 75, 63, 62,
  75, 76, 64, 63,
  76, 77, 65, 64,
  77, 78, 66, 65,
  78, 79, 67, 66,
  79, 80, 68, 67,
  80, 81, 69, 68,
  81, 82, 70, 69,
  82, 83, 71, 70,
  83, 84, 72, 71,
  84, 217, 205, 72,
  85, 86, 74, 73,
  86, 87, 75, 74,
  87, 88, 76, 75,
  88, 89, 77, 76,
  89, 90, 78, 77,
  90, 91, 79, 78,
  91, 92, 80, 79,
  92, 93, 81, 80,
  93, 94, 82, 81,
  94, 95, 83, 82,
  95, 96, 84, 83,
  96, 229, 217, 84,
  97, 98, 86, 85,
  98, 99, 87, 86,
  99, 100, 88, 87,
  100, 101, 89, 88,
  101, 102, 90, 89,
  102, 103, 91, 90,
  103, 104, 92, 91,
  104, 105, 93, 92,
  105, 106, 94, 93,
  106, 107, 95, 94,
  107, 108, 96, 95,
  108, 241, 229, 96,
  109, 110, 98, 97,
  110, 111, 99, 98,
  111, 112, 100, 99,
  112, 113, 101, 100,
  113, 114, 102, 101,
  114, 115, 103, 102,
  115, 116, 104, 103,
  116, 117, 105, 104,
  117, 118, 106, 105,
  118, 119, 107, 106,
  119, 120, 108, 107,
  120, 253, 241, 108,
  121, 122, 110, 109,
  122, 123, 111, 110,
  123, 124, 112, 111,
  124, 125, 113, 112,
  125, 126, 114, 113,
  126, 127, 115, 114,
  127, 128, 116, 115,
  128, 129, 117, 116,
  129, 130, 118, 117,
  130, 131, 119, 118,
  131, 132, 120, 119,
  132, 265, 253, 120,
  133, 134, 122, 121,
  134, 135, 123, 122,
  135, 136, 124, 123,
  136, 137, 125, 124,
  137, 138, 126, 125,
  138, 139, 127, 126,
  139, 140, 128, 127,
  140, 141, 129, 128,
  141, 142, 130, 129,
  142, 143, 131, 130,
  143, 144, 132, 131,
  144, 277, 265, 132,
  842, 830, 134, 133,
  830, 818, 135, 134,
  818, 806, 136, 135,
  806, 794, 137, 136,
  794, 782, 138, 137,
  782, 770, 139, 138,
  770, 758, 140, 139,
  758, 746, 141, 140,
  746, 734, 142, 141,
  734, 722, 143, 142,
  722, 710, 144, 143,
  710, 698, 277, 144,
  157, 158, 146, 145,
  158, 159, 147, 146,
  159, 160, 148, 147,
  160, 161, 149, 148,
  161, 162, 150, 149,
  162, 163, 151, 150,
  163, 164, 152, 151,
  164, 165, 153, 152,
  165, 166, 154, 153,
  166, 167, 155, 154,
  167, 168, 156, 155,
  168, 301, 289, 156,
  169, 170, 158, 157,
  170, 171, 159, 158,
  171, 172, 160, 159,
  172, 173, 161, 160,
  173, 174, 162, 161,
  174, 175, 163, 162,
  175, 176, 164, 163,
  176, 177, 165, 164,
  177, 178, 166, 165,
  178, 179, 167, 166,
  179, 180, 168, 167,
  180, 313, 301, 168,
  181, 182, 170, 169,
  182, 183, 171, 170,
  183, 184, 172, 171,
  184, 185, 173, 172,
  185, 186, 174, 173,
  186, 187, 175, 174,
  187, 188, 176, 175,
  188, 189, 177, 176,
  189, 190, 178, 177,
  190, 191, 179, 178,
  191, 192, 180, 179,
  192, 325, 313, 180,
  193, 194, 182, 181,
  194, 195, 183, 182,
  195, 196, 184, 183,
  196, 197, 185, 184,
  197, 198, 186, 185,
  198, 199, 187, 186,
  199, 200, 188, 187,
  200, 201, 189, 188,
  201, 202, 190, 189,
  202, 203, 191, 190,
  203, 204, 192, 191,
  204, 337, 325, 192,
  205, 206, 194, 193,
  206, 207, 195, 194,
  207, 208, 196, 195,
  208, 209, 197, 196,
  209, 210, 198, 197,
  210, 211, 199, 198,
  211, 212, 200, 199,
  212, 213, 201, 200,
  213, 214, 202, 201,
  214, 215, 203, 202,
  215, 216, 204, 203,
  216, 349, 337, 204,
  217, 218, 206, 205,
  218, 219, 207, 206,
  219, 220, 208, 207,
  220, 221, 209, 208,
  221, 222, 210, 209,
  222, 223, 211, 210,
  223, 224, 212, 211,
  224, 225, 213, 212,
  225, 226, 214, 213,
  226, 227, 215, 214,
  227, 228, 216, 215,
  228, 361, 349, 216,
  229, 230, 218, 217,
  230, 231, 219, 218,
  231, 232, 220, 219,
  232, 233, 221, 220,
  233, 234, 222, 221,
  234, 235, 223, 222,
  235, 236, 224, 223,
  236, 237, 225, 224,
  237, 238, 226, 225,
  238, 239, 227, 226,
  239, 240, 228, 227,
  240, 373, 361, 228,
  241, 242, 230, 229,
  242, 243, 231, 230,
  243, 244, 232, 231,
  244, 245, 233, 232,
  245, 246, 234, 233,
  246, 247, 235, 234,
  247, 248, 236, 235,
  248, 249, 237, 236,
  249, 250, 238, 237,
  250, 251, 239, 238,
  251, 252, 240, 239,
  252, 385, 373, 240,
  253, 254, 242, 241,
  254, 255, 243, 242,
  255, 256, 244, 243,
  256, 257, 245, 244,
  257, 258, 246, 245,
  258, 259, 247, 246,
  259, 260, 248, 247,
  260, 261, 249, 248,
  261, 262, 250, 249,
  262, 263, 251, 250,
  263, 264, 252, 251,
  264, 397, 385, 252,
  265, 266, 254, 253,
  266, 267, 255, 254,
  267, 268, 256, 255,
  268, 269, 257, 256,
  269, 270, 258, 257,
  270, 271, 259, 258,
  271, 272, 260, 259,
  272, 273, 261, 260,
  273, 274, 262, 261,
  274, 275, 263, 262,
  275, 276, 264, 263,
  276, 409, 397, 264,
  277, 278, 266, 265,
  278, 279, 267, 266,
  279, 280, 268, 267,
  280, 281, 269, 268,
  281, 282, 270, 269,
  282, 283, 271, 270,
  283, 284, 272, 271,
  284, 285, 273, 272,
  285, 286, 274, 273,
  286, 287, 275, 274,
  287, 288, 276, 275,
  288, 421, 409, 276,
  698, 699, 278, 277,
  699, 700, 279, 278,
  700, 701, 280, 279,
  701, 702, 281, 280,
  702, 703, 282, 281,
  703, 704, 283, 282,
  704, 705, 284, 283,
  705, 706, 285, 284,
  706, 707, 286, 285,
  707, 708, 287, 286,
  708, 709, 288, 287,
  709, 854, 421, 288,
  302, 290, 289, 301,
  303, 291, 290, 302,
  304, 292, 291, 303,
  305, 293, 292, 304,
  306, 294, 293, 305,
  307, 295, 294, 306,
  308, 296, 295, 307,
  309, 297, 296, 308,
  310, 298, 297, 309,
  311, 299, 298, 310,
  312, 300, 299, 311,
  445, 433, 300, 312,
  314, 302, 301, 313,
  315, 303, 302, 314,
  316, 304, 303, 315,
  317, 305, 304, 316,
  318, 306, 305, 317,
  319, 307, 306, 318,
  320, 308, 307, 319,
  321, 309, 308, 320,
  322, 310, 309, 321,
  323, 311, 310, 322,
  324, 312, 311, 323,
  457, 445, 312, 324,
  326, 314, 313, 325,
  327, 315, 314, 326,
  328, 316, 315, 327,
  329, 317, 316, 328,
  330, 318, 317, 329,
  331, 319, 318, 330,
  332, 320, 319, 331,
  333, 321, 320, 332,
  334, 322, 321, 333,
  335, 323, 322, 334,
  336, 324, 323, 335,
  469, 457, 324, 336,
  338, 326, 325, 337,
  339, 327, 326, 338,
  340, 328, 327, 339,
  341, 329, 328, 340,
  342, 330, 329, 341,
  343, 331, 330, 342,
  344, 332, 331, 343,
  345, 333, 332, 344,
  346, 334, 333, 345,
  347, 335, 334, 346,
  348, 336, 335, 347,
  481, 469, 336, 348,
  350, 338, 337, 349,
  351, 339, 338, 350,
  352, 340, 339, 351,
  353, 341, 340, 352,
  354, 342, 341, 353,
  355, 343, 342, 354,
  356, 344, 343, 355,
  357, 345, 344, 356,
  358, 346, 345, 357,
  359, 347, 346, 358,
  360, 348, 347, 359,
  493, 481, 348, 360,
  362, 350, 349, 361,
  363, 351, 350, 362,
  364, 352, 351, 363,
  365, 353, 352, 364,
  366, 354, 353, 365,
  367, 355, 354, 366,
  368, 356, 355, 367,
  369, 357, 356, 368,
  370, 358, 357, 369,
  371, 359, 358, 370,
  372, 360, 359, 371,
  505, 493, 360, 372,
  374, 362, 361, 373,
  375, 363, 362, 374,
  376, 364, 363, 375,
  377, 365, 364, 376,
  378, 366, 365, 377,
  379, 367, 366, 378,
  380, 368, 367, 379,
  381, 369, 368, 380,
  382, 370, 369, 381,
  383, 371, 370, 382,
  384, 372, 371, 383,
  517, 505, 372, 384,
  386, 374, 373, 385,
  387, 375, 374, 386,
  388, 376, 375, 387,
  389, 377, 376, 388,
  390, 378, 377, 389,
  391, 379, 378, 390,
  392, 380, 379, 391,
  393, 381, 380, 392,
  394, 382, 381, 393,
  395, 383, 382, 394,
  396, 384, 383, 395,
  529, 517, 384, 396,
  398, 386, 385, 397,
  399, 387, 386, 398,
  400, 388, 387, 399,
  401, 389, 388, 400,
  402, 390, 389, 401,
  403, 391, 390, 402,
  404, 392, 391, 403,
  405, 393, 392, 404,
  406, 394, 393, 405,
  407, 395, 394, 406,
  408, 396, 395, 407,
  541, 529, 396, 408,
  410, 398, 397, 409,
  411, 399, 398, 410,
  412, 400, 399, 411,
  413, 401, 400, 412,
  414, 402, 401, 413,
  415, 403, 402, 414,
  416, 404, 403, 415,
  417, 405, 404, 416,
  418, 406, 405, 417,
  419, 407, 406, 418,
  420, 408, 407, 419,
  553, 541, 408, 420,
  422, 410, 409, 421,
  423, 411, 410, 422,
  424, 412, 411, 423,
  425, 413, 412, 424,
  426, 414, 413, 425,
  427, 415, 414, 426,
  428, 416, 415, 427,
  429, 417, 416, 428,
  430, 418, 417, 429,
  431, 419, 418, 430,
  432, 420, 419, 431,
  565, 553, 420, 432,
  855, 422, 421, 854,
  856, 423, 422, 855,
  857, 424, 423, 856,
  858, 425, 424, 857,
  859, 426, 425, 858,
  860, 427, 426, 859,
  861, 428, 427, 860,
  862, 429, 428, 861,
  863, 430, 429, 862,
  864, 431, 430, 863,
  865, 432, 431, 864,
  866, 565, 432, 865,
  446, 434, 433, 445,
  447, 435, 434, 446,
  448, 436, 435, 447,
  449, 437, 436, 448,
  450, 438, 437, 449,
  451, 439, 438, 450,
  452, 440, 439, 451,
  453, 441, 440, 452,
  454, 442, 441, 453,
  455, 443, 442, 454,
  456, 444, 443, 455,
  13, 1, 444, 456,
  458, 446, 445, 457,
  459, 447, 446, 458,
  460, 448, 447, 459,
  461, 449, 448, 460,
  462, 450, 449, 461,
  463, 451, 450, 462,
  464, 452, 451, 463,
  465, 453, 452, 464,
  466, 454, 453, 465,
  467, 455, 454, 466,
  468, 456, 455, 467,
  25, 13, 456, 468,
  470, 458, 457, 469,
  471, 459, 458, 470,
  472, 460, 459, 471,
  473, 461, 460, 472,
  474, 462, 461, 473,
  475, 463, 462, 474,
  476, 464, 463, 475,
  477, 465, 464, 476,
  478, 466, 465, 477,
  479, 467, 466, 478,
  480, 468, 467, 479,
  37, 25, 468, 480,
  482, 470, 469, 481,
  483, 471, 470, 482,
  484, 472, 471, 483,
  485, 473, 472, 484,
  486, 474, 473, 485,
  487, 475, 474, 486,
  488, 476, 475, 487,
  489, 477, 476, 488,
  490, 478, 477, 489,
  491, 479, 478, 490,
  492, 480, 479, 491,
  49, 37, 480, 492,
  494, 482, 481, 493,
  495, 483, 482, 494,
  496, 484, 483, 495,
  497, 485, 484, 496,
  498, 486, 485, 497,
  499, 487, 486, 498,
  500, 488, 487, 499,
  501, 489, 488, 500,
  502, 490, 489, 501,
  503, 491, 490, 502,
  504, 492, 491, 503,
  61, 49, 492, 504,
  506, 494, 493, 505,
  507, 495, 494, 506,
  508, 496, 495, 507,
  509, 497, 496, 508,
  510, 498, 497, 509,
  511, 499, 498, 510,
  512, 500, 499, 511,
  513, 501, 500, 512,
  514, 502, 501, 513,
  515, 503, 502, 514,
  516, 504, 503, 515,
  73, 61, 504, 516,
  518, 506, 505, 517,
  519, 507, 506, 518,
  520, 508, 507, 519,
  521, 509, 508, 520,
  522, 510, 509, 521,
  523, 511, 510, 522,
  524, 512, 511, 523,
  525, 513, 512, 524,
  526, 514, 513, 525,
  527, 515, 514, 526,
  528, 516, 515, 527,
  85, 73, 516, 528,
  530, 518, 517, 529,
  531, 519, 518, 530,
  532, 520, 519, 531,
  533, 521, 520, 532,
  534, 522, 521, 533,
  535, 523, 522, 534,
  536, 524, 523, 535,
  537, 525, 524, 536,
  538, 526, 525, 537,
  539, 527, 526, 538,
  540, 528, 527, 539,
  97, 85, 528, 540,
  542, 530, 529, 541,
  543, 531, 530, 542,
  544, 532, 531, 543,
  545, 533, 532, 544,
  546, 534, 533, 545,
  547, 535, 534, 546,
  548, 536, 535, 547,
  549, 537, 536, 548,
  550, 538, 537, 549,
  551, 539, 538, 550,
  552, 540, 539, 551,
  109, 97, 540, 552,
  554, 542, 541, 553,
  555, 543, 542, 554,
  556, 544, 543, 555,
  557, 545, 544, 556,
  558, 546, 545, 557,
  559, 547, 546, 558,
  560, 548, 547, 559,
  561, 549, 548, 560,
  562, 550, 549, 561,
  563, 551, 550, 562,
  564, 552, 551, 563,
  121, 109, 552, 564,
  566, 554, 553, 565,
  567, 555, 554, 566,
  568, 556, 555, 567,
  569, 557, 556, 568,
  570, 558, 557, 569,
  571, 559, 558, 570,
  572, 560, 559, 571,
  573, 561, 560, 572,
  574, 562, 561, 573,
  575, 563, 562, 574,
  576, 564, 563, 575,
  133, 121, 564, 576,
  853, 566, 565, 866,
  852, 567, 566, 853,
  851, 568, 567, 852,
  850, 569, 568, 851,
  849, 570, 569, 850,
  848, 571, 570, 849,
  847, 572, 571, 848,
  846, 573, 572, 847,
  845, 574, 573, 846,
  844, 575, 574, 845,
  843, 576, 575, 844,
  842, 133, 576, 843,
  1, 2, 577, 444,
  444, 577, 578, 443,
  443, 578, 579, 442,
  442, 579, 580, 441,
  441, 580, 581, 440,
  440, 581, 582, 439,
  439, 582, 583, 438,
  438, 583, 584, 437,
  437, 584, 585, 436,
  436, 585, 586, 435,
  435, 586, 587, 434,
  434, 587, 300, 433,
  2, 3, 588, 577,
  577, 588, 589, 578,
  578, 589, 590, 579,
  579, 590, 591, 580,
  580, 591, 592, 581,
  581, 592, 593, 582,
  582, 593, 594, 583,
  583, 594, 595, 584,
  584, 595, 596, 585,
  585, 596, 597, 586,
  586, 597, 598, 587,
  587, 598, 299, 300,
  3, 4, 599, 588,
  588, 599, 600, 589,
  589, 600, 601, 590,
  590, 601, 602, 591,
  591, 602, 603, 592,
  592, 603, 604, 593,
  593, 604, 605, 594,
  594, 605, 606, 595,
  595, 606, 607, 596,
  596, 607, 608, 597,
  597, 608, 609, 598,
  598, 609, 298, 299,
  4, 5, 610, 599,
  599, 610, 611, 600,
  600, 611, 612, 601,
  601, 612, 613, 602,
  602, 613, 614, 603,
  603, 614, 615, 604,
  604, 615, 616, 605,
  605, 616, 617, 606,
  606, 617, 618, 607,
  607, 618, 619, 608,
  608, 619, 620, 609,
  609, 620, 297, 298,
  5, 6, 621, 610,
  610, 621, 622, 611,
  611, 622, 623, 612,
  612, 623, 624, 613,
  613, 624, 625, 614,
  614, 625, 626, 615,
  615, 626, 627, 616,
  616, 627, 628, 617,
  617, 628, 629, 618,
  618, 629, 630, 619,
  619, 630, 631, 620,
  620, 631, 296, 297,
  6, 7, 632, 621,
  621, 632, 633, 622,
  622, 633, 634, 623,
  623, 634, 635, 624,
  624, 635, 636, 625,
  625, 636, 637, 626,
  626, 637, 638, 627,
  627, 638, 639, 628,
  628, 639, 640, 629,
  629, 640, 641, 630,
  630, 641, 642, 631,
  631, 642, 295, 296,
  7, 8, 643, 632,
  632, 643, 644, 633,
  633, 644, 645, 634,
  634, 645, 646, 635,
  635, 646, 647, 636,
  636, 647, 648, 637,
  637, 648, 649, 638,
  638, 649, 650, 639,
  639, 650, 651, 640,
  640, 651, 652, 641,
  641, 652, 653, 642,
  642, 653, 294, 295,
  8, 9, 654, 643,
  643, 654, 655, 644,
  644, 655, 656, 645,
  645, 656, 657, 646,
  646, 657, 658, 647,
  647, 658, 659, 648,
  648, 659, 660, 649,
  649, 660, 661, 650,
  650, 661, 662, 651,
  651, 662, 663, 652,
  652, 663, 664, 653,
  653, 664, 293, 294,
  9, 10, 665, 654,
  654, 665, 666, 655,
  655, 666, 667, 656,
  656, 667, 668, 657,
  657, 668, 669, 658,
  658, 669, 670, 659,
  659, 670, 671, 660,
  660, 671, 672, 661,
  661, 672, 673, 662,
  662, 673, 674, 663,
  663, 674, 675, 664,
  664, 675, 292, 293,
  10, 11, 676, 665,
  665, 676, 677, 666,
  666, 677, 678, 667,
  667, 678, 679, 668,
  668, 679, 680, 669,
  669, 680, 681, 670,
  670, 681, 682, 671,
  671, 682, 683, 672,
  672, 683, 684, 673,
  673, 684, 685, 674,
  674, 685, 686, 675,
  675, 686, 291, 292,
  11, 12, 687, 676,
  676, 687, 688, 677,
  677, 688, 689, 678,
  678, 689, 690, 679,
  679, 690, 691, 680,
  680, 691, 692, 681,
  681, 692, 693, 682,
  682, 693, 694, 683,
  683, 694, 695, 684,
  684, 695, 696, 685,
  685, 696, 697, 686,
  686, 697, 290, 291,
  12, 145, 146, 687,
  687, 146, 147, 688,
  688, 147, 148, 689,
  689, 148, 149, 690,
  690, 149, 150, 691,
  691, 150, 151, 692,
  692, 151, 152, 693,
  693, 152, 153, 694,
  694, 153, 154, 695,
  695, 154, 155, 696,
  696, 155, 156, 697,
  697, 156, 289, 290,
  710, 711, 699, 698,
  711, 712, 700, 699,
  712, 713, 701, 700,
  713, 714, 702, 701,
  714, 715, 703, 702,
  715, 716, 704, 703,
  716, 717, 705, 704,
  717, 718, 706, 705,
  718, 719, 707, 706,
  719, 720, 708, 707,
  720, 721, 709, 708,
  721, 855, 854, 709,
  722, 723, 711, 710,
  723, 724, 712, 711,
  724, 725, 713, 712,
  725, 726, 714, 713,
  726, 727, 715, 714,
  727, 728, 716, 715,
  728, 729, 717, 716,
  729, 730, 718, 717,
  730, 731, 719, 718,
  731, 732, 720, 719,
  732, 733, 721, 720,
  733, 856, 855, 721,
  734, 735, 723, 722,
  735, 736, 724, 723,
  736, 737, 725, 724,
  737, 738, 726, 725,
  738, 739, 727, 726,
  739, 740, 728, 727,
  740, 741, 729, 728,
  741, 742, 730, 729,
  742, 743, 731, 730,
  743, 744, 732, 731,
  744, 745, 733, 732,
  745, 857, 856, 733,
  746, 747, 735, 734,
  747, 748, 736, 735,
  748, 749, 737, 736,
  749, 750, 738, 737,
  750, 751, 739, 738,
  751, 752, 740, 739,
  752, 753, 741, 740,
  753, 754, 742, 741,
  754, 755, 743, 742,
  755, 756, 744, 743,
  756, 757, 745, 744,
  757, 858, 857, 745,
  758, 759, 747, 746,
  759, 760, 748, 747,
  760, 761, 749, 748,
  761, 762, 750, 749,
  762, 763, 751, 750,
  763, 764, 752, 751,
  764, 765, 753, 752,
  765, 766, 754, 753,
  766, 767, 755, 754,
  767, 768, 756, 755,
  768, 769, 757, 756,
  769, 859, 858, 757,
  770, 771, 759, 758,
  771, 772, 760, 759,
  772, 773, 761, 760,
  773, 774, 762, 761,
  774, 775, 763, 762,
  775, 776, 764, 763,
  776, 777, 765, 764,
  777, 778, 766, 765,
  778, 779, 767, 766,
  779, 780, 768, 767,
  780, 781, 769, 768,
  781, 860, 859, 769,
  782, 783, 771, 770,
  783, 784, 772, 771,
  784, 785, 773, 772,
  785, 786, 774, 773,
  786, 787, 775, 774,
  787, 788, 776, 775,
  788, 789, 777, 776,
  789, 790, 778, 777,
  790, 791, 779, 778,
  791, 792, 780, 779,
  792, 793, 781, 780,
  793, 861, 860, 781,
  794, 795, 783, 782,
  795, 796, 784, 783,
  796, 797, 785, 784,
  797, 798, 786, 785,
  798, 799, 787, 786,
  799, 800, 788, 787,
  800, 801, 789, 788,
  801, 802, 790, 789,
  802, 803, 791, 790,
  803, 804, 792, 791,
  804, 805, 793, 792,
  805, 862, 861, 793,
  806, 807, 795, 794,
  807, 808, 796, 795,
  808, 809, 797, 796,
  809, 810, 798, 797,
  810, 811, 799, 798,
  811, 812, 800, 799,
  812, 813, 801, 800,
  813, 814, 802, 801,
  814, 815, 803, 802,
  815, 816, 804, 803,
  816, 817, 805, 804,
  817, 863, 862, 805,
  818, 819, 807, 806,
  819, 820, 808, 807,
  820, 821, 809, 808,
  821, 822, 810, 809,
  822, 823, 811, 810,
  823, 824, 812, 811,
  824, 825, 813, 812,
  825, 826, 814, 813,
  826, 827, 815, 814,
  827, 828, 816, 815,
  828, 829, 817, 816,
  829, 864, 863, 817,
  830, 831, 819, 818,
  831, 832, 820, 819,
  832, 833, 821, 820,
  833, 834, 822, 821,
  834, 835, 823, 822,
  835, 836, 824, 823,
  836, 837, 825, 824,
  837, 838, 826, 825,
  838, 839, 827, 826,
  839, 840, 828, 827,
  840, 841, 829, 828,
  841, 865, 864, 829,
  842, 843, 831, 830,
  843, 844, 832, 831,
  844, 845, 833, 832,
  845, 846, 834, 833,
  846, 847, 835, 834,
  847, 848, 836, 835,
  848, 849, 837, 836,
  849, 850, 838, 837,
  850, 851, 839, 838,
  851, 852, 840, 839,
  852, 853, 841, 840,
  853, 866, 865, 841 ;

 dynamics_edge_nodes =
  1, 2,
  13, 1,
  14, 13,
  2, 3,
  14, 2,
  15, 14,
  3, 4,
  15, 3,
  16, 15,
  4, 5,
  16, 4,
  17, 16,
  5, 6,
  17, 5,
  18, 17,
  6, 7,
  18, 6,
  19, 18,
  7, 8,
  19, 7,
  20, 19,
  8, 9,
  20, 8,
  21, 20,
  9, 10,
  21, 9,
  22, 21,
  10, 11,
  22, 10,
  23, 22,
  11, 12,
  23, 11,
  24, 23,
  12, 145,
  24, 12,
  157, 24,
  25, 13,
  26, 25,
  26, 14,
  27, 26,
  27, 15,
  28, 27,
  28, 16,
  29, 28,
  29, 17,
  30, 29,
  30, 18,
  31, 30,
  31, 19,
  32, 31,
  32, 20,
  33, 32,
  33, 21,
  34, 33,
  34, 22,
  35, 34,
  35, 23,
  36, 35,
  36, 24,
  169, 36,
  37, 25,
  38, 37,
  38, 26,
  39, 38,
  39, 27,
  40, 39,
  40, 28,
  41, 40,
  41, 29,
  42, 41,
  42, 30,
  43, 42,
  43, 31,
  44, 43,
  44, 32,
  45, 44,
  45, 33,
  46, 45,
  46, 34,
  47, 46,
  47, 35,
  48, 47,
  48, 36,
  181, 48,
  49, 37,
  50, 49,
  50, 38,
  51, 50,
  51, 39,
  52, 51,
  52, 40,
  53, 52,
  53, 41,
  54, 53,
  54, 42,
  55, 54,
  55, 43,
  56, 55,
  56, 44,
  57, 56,
  57, 45,
  58, 57,
  58, 46,
  59, 58,
  59, 47,
  60, 59,
  60, 48,
  193, 60,
  61, 49,
  62, 61,
  62, 50,
  63, 62,
  63, 51,
  64, 63,
  64, 52,
  65, 64,
  65, 53,
  66, 65,
  66, 54,
  67, 66,
  67, 55,
  68, 67,
  68, 56,
  69, 68,
  69, 57,
  70, 69,
  70, 58,
  71, 70,
  71, 59,
  72, 71,
  72, 60,
  205, 72,
  73, 61,
  74, 73,
  74, 62,
  75, 74,
  75, 63,
  76, 75,
  76, 64,
  77, 76,
  77, 65,
  78, 77,
  78, 66,
  79, 78,
  79, 67,
  80, 79,
  80, 68,
  81, 80,
  81, 69,
  82, 81,
  82, 70,
  83, 82,
  83, 71,
  84, 83,
  84, 72,
  217, 84,
  85, 73,
  86, 85,
  86, 74,
  87, 86,
  87, 75,
  88, 87,
  88, 76,
  89, 88,
  89, 77,
  90, 89,
  90, 78,
  91, 90,
  91, 79,
  92, 91,
  92, 80,
  93, 92,
  93, 81,
  94, 93,
  94, 82,
  95, 94,
  95, 83,
  96, 95,
  96, 84,
  229, 96,
  97, 85,
  98, 97,
  98, 86,
  99, 98,
  99, 87,
  100, 99,
  100, 88,
  101, 100,
  101, 89,
  102, 101,
  102, 90,
  103, 102,
  103, 91,
  104, 103,
  104, 92,
  105, 104,
  105, 93,
  106, 105,
  106, 94,
  107, 106,
  107, 95,
  108, 107,
  108, 96,
  241, 108,
  109, 97,
  110, 109,
  110, 98,
  111, 110,
  111, 99,
  112, 111,
  112, 100,
  113, 112,
  113, 101,
  114, 113,
  114, 102,
  115, 114,
  115, 103,
  116, 115,
  116, 104,
  117, 116,
  117, 105,
  118, 117,
  118, 106,
  119, 118,
  119, 107,
  120, 119,
  120, 108,
  253, 120,
  121, 109,
  122, 121,
  122, 110,
  123, 122,
  123, 111,
  124, 123,
  124, 112,
  125, 124,
  125, 113,
  126, 125,
  126, 114,
  127, 126,
  127, 115,
  128, 127,
  128, 116,
  129, 128,
  129, 117,
  130, 129,
  130, 118,
  131, 130,
  131, 119,
  132, 131,
  132, 120,
  265, 132,
  133, 121,
  134, 133,
  134, 122,
  135, 134,
  135, 123,
  136, 135,
  136, 124,
  137, 136,
  137, 125,
  138, 137,
  138, 126,
  139, 138,
  139, 127,
  140, 139,
  140, 128,
  141, 140,
  141, 129,
  142, 141,
  142, 130,
  143, 142,
  143, 131,
  144, 143,
  144, 132,
  277, 144,
  842, 133,
  830, 842,
  830, 134,
  818, 830,
  818, 135,
  806, 818,
  806, 136,
  794, 806,
  794, 137,
  782, 794,
  782, 138,
  770, 782,
  770, 139,
  758, 770,
  758, 140,
  746, 758,
  746, 141,
  734, 746,
  734, 142,
  722, 734,
  722, 143,
  710, 722,
  710, 144,
  698, 710,
  145, 146,
  157, 145,
  158, 157,
  146, 147,
  158, 146,
  159, 158,
  147, 148,
  159, 147,
  160, 159,
  148, 149,
  160, 148,
  161, 160,
  149, 150,
  161, 149,
  162, 161,
  150, 151,
  162, 150,
  163, 162,
  151, 152,
  163, 151,
  164, 163,
  152, 153,
  164, 152,
  165, 164,
  153, 154,
  165, 153,
  166, 165,
  154, 155,
  166, 154,
  167, 166,
  155, 156,
  167, 155,
  168, 167,
  156, 289,
  168, 156,
  301, 168,
  169, 157,
  170, 169,
  170, 158,
  171, 170,
  171, 159,
  172, 171,
  172, 160,
  173, 172,
  173, 161,
  174, 173,
  174, 162,
  175, 174,
  175, 163,
  176, 175,
  176, 164,
  177, 176,
  177, 165,
  178, 177,
  178, 166,
  179, 178,
  179, 167,
  180, 179,
  180, 168,
  313, 180,
  181, 169,
  182, 181,
  182, 170,
  183, 182,
  183, 171,
  184, 183,
  184, 172,
  185, 184,
  185, 173,
  186, 185,
  186, 174,
  187, 186,
  187, 175,
  188, 187,
  188, 176,
  189, 188,
  189, 177,
  190, 189,
  190, 178,
  191, 190,
  191, 179,
  192, 191,
  192, 180,
  325, 192,
  193, 181,
  194, 193,
  194, 182,
  195, 194,
  195, 183,
  196, 195,
  196, 184,
  197, 196,
  197, 185,
  198, 197,
  198, 186,
  199, 198,
  199, 187,
  200, 199,
  200, 188,
  201, 200,
  201, 189,
  202, 201,
  202, 190,
  203, 202,
  203, 191,
  204, 203,
  204, 192,
  337, 204,
  205, 193,
  206, 205,
  206, 194,
  207, 206,
  207, 195,
  208, 207,
  208, 196,
  209, 208,
  209, 197,
  210, 209,
  210, 198,
  211, 210,
  211, 199,
  212, 211,
  212, 200,
  213, 212,
  213, 201,
  214, 213,
  214, 202,
  215, 214,
  215, 203,
  216, 215,
  216, 204,
  349, 216,
  217, 205,
  218, 217,
  218, 206,
  219, 218,
  219, 207,
  220, 219,
  220, 208,
  221, 220,
  221, 209,
  222, 221,
  222, 210,
  223, 222,
  223, 211,
  224, 223,
  224, 212,
  225, 224,
  225, 213,
  226, 225,
  226, 214,
  227, 226,
  227, 215,
  228, 227,
  228, 216,
  361, 228,
  229, 217,
  230, 229,
  230, 218,
  231, 230,
  231, 219,
  232, 231,
  232, 220,
  233, 232,
  233, 221,
  234, 233,
  234, 222,
  235, 234,
  235, 223,
  236, 235,
  236, 224,
  237, 236,
  237, 225,
  238, 237,
  238, 226,
  239, 238,
  239, 227,
  240, 239,
  240, 228,
  373, 240,
  241, 229,
  242, 241,
  242, 230,
  243, 242,
  243, 231,
  244, 243,
  244, 232,
  245, 244,
  245, 233,
  246, 245,
  246, 234,
  247, 246,
  247, 235,
  248, 247,
  248, 236,
  249, 248,
  249, 237,
  250, 249,
  250, 238,
  251, 250,
  251, 239,
  252, 251,
  252, 240,
  385, 252,
  253, 241,
  254, 253,
  254, 242,
  255, 254,
  255, 243,
  256, 255,
  256, 244,
  257, 256,
  257, 245,
  258, 257,
  258, 246,
  259, 258,
  259, 247,
  260, 259,
  260, 248,
  261, 260,
  261, 249,
  262, 261,
  262, 250,
  263, 262,
  263, 251,
  264, 263,
  264, 252,
  397, 264,
  265, 253,
  266, 265,
  266, 254,
  267, 266,
  267, 255,
  268, 267,
  268, 256,
  269, 268,
  269, 257,
  270, 269,
  270, 258,
  271, 270,
  271, 259,
  272, 271,
  272, 260,
  273, 272,
  273, 261,
  274, 273,
  274, 262,
  275, 274,
  275, 263,
  276, 275,
  276, 264,
  409, 276,
  277, 265,
  278, 277,
  278, 266,
  279, 278,
  279, 267,
  280, 279,
  280, 268,
  281, 280,
  281, 269,
  282, 281,
  282, 270,
  283, 282,
  283, 271,
  284, 283,
  284, 272,
  285, 284,
  285, 273,
  286, 285,
  286, 274,
  287, 286,
  287, 275,
  288, 287,
  288, 276,
  421, 288,
  698, 277,
  699, 698,
  699, 278,
  700, 699,
  700, 279,
  701, 700,
  701, 280,
  702, 701,
  702, 281,
  703, 702,
  703, 282,
  704, 703,
  704, 283,
  705, 704,
  705, 284,
  706, 705,
  706, 285,
  707, 706,
  707, 286,
  708, 707,
  708, 287,
  709, 708,
  709, 288,
  854, 709,
  289, 290,
  301, 289,
  302, 301,
  290, 291,
  302, 290,
  303, 302,
  291, 292,
  303, 291,
  304, 303,
  292, 293,
  304, 292,
  305, 304,
  293, 294,
  305, 293,
  306, 305,
  294, 295,
  306, 294,
  307, 306,
  295, 296,
  307, 295,
  308, 307,
  296, 297,
  308, 296,
  309, 308,
  297, 298,
  309, 297,
  310, 309,
  298, 299,
  310, 298,
  311, 310,
  299, 300,
  311, 299,
  312, 311,
  300, 433,
  312, 300,
  445, 312,
  313, 301,
  314, 313,
  314, 302,
  315, 314,
  315, 303,
  316, 315,
  316, 304,
  317, 316,
  317, 305,
  318, 317,
  318, 306,
  319, 318,
  319, 307,
  320, 319,
  320, 308,
  321, 320,
  321, 309,
  322, 321,
  322, 310,
  323, 322,
  323, 311,
  324, 323,
  324, 312,
  457, 324,
  325, 313,
  326, 325,
  326, 314,
  327, 326,
  327, 315,
  328, 327,
  328, 316,
  329, 328,
  329, 317,
  330, 329,
  330, 318,
  331, 330,
  331, 319,
  332, 331,
  332, 320,
  333, 332,
  333, 321,
  334, 333,
  334, 322,
  335, 334,
  335, 323,
  336, 335,
  336, 324,
  469, 336,
  337, 325,
  338, 337,
  338, 326,
  339, 338,
  339, 327,
  340, 339,
  340, 328,
  341, 340,
  341, 329,
  342, 341,
  342, 330,
  343, 342,
  343, 331,
  344, 343,
  344, 332,
  345, 344,
  345, 333,
  346, 345,
  346, 334,
  347, 346,
  347, 335,
  348, 347,
  348, 336,
  481, 348,
  349, 337,
  350, 349,
  350, 338,
  351, 350,
  351, 339,
  352, 351,
  352, 340,
  353, 352,
  353, 341,
  354, 353,
  354, 342,
  355, 354,
  355, 343,
  356, 355,
  356, 344,
  357, 356,
  357, 345,
  358, 357,
  358, 346,
  359, 358,
  359, 347,
  360, 359,
  360, 348,
  493, 360,
  361, 349,
  362, 361,
  362, 350,
  363, 362,
  363, 351,
  364, 363,
  364, 352,
  365, 364,
  365, 353,
  366, 365,
  366, 354,
  367, 366,
  367, 355,
  368, 367,
  368, 356,
  369, 368,
  369, 357,
  370, 369,
  370, 358,
  371, 370,
  371, 359,
  372, 371,
  372, 360,
  505, 372,
  373, 361,
  374, 373,
  374, 362,
  375, 374,
  375, 363,
  376, 375,
  376, 364,
  377, 376,
  377, 365,
  378, 377,
  378, 366,
  379, 378,
  379, 367,
  380, 379,
  380, 368,
  381, 380,
  381, 369,
  382, 381,
  382, 370,
  383, 382,
  383, 371,
  384, 383,
  384, 372,
  517, 384,
  385, 373,
  386, 385,
  386, 374,
  387, 386,
  387, 375,
  388, 387,
  388, 376,
  389, 388,
  389, 377,
  390, 389,
  390, 378,
  391, 390,
  391, 379,
  392, 391,
  392, 380,
  393, 392,
  393, 381,
  394, 393,
  394, 382,
  395, 394,
  395, 383,
  396, 395,
  396, 384,
  529, 396,
  397, 385,
  398, 397,
  398, 386,
  399, 398,
  399, 387,
  400, 399,
  400, 388,
  401, 400,
  401, 389,
  402, 401,
  402, 390,
  403, 402,
  403, 391,
  404, 403,
  404, 392,
  405, 404,
  405, 393,
  406, 405,
  406, 394,
  407, 406,
  407, 395,
  408, 407,
  408, 396,
  541, 408,
  409, 397,
  410, 409,
  410, 398,
  411, 410,
  411, 399,
  412, 411,
  412, 400,
  413, 412,
  413, 401,
  414, 413,
  414, 402,
  415, 414,
  415, 403,
  416, 415,
  416, 404,
  417, 416,
  417, 405,
  418, 417,
  418, 406,
  419, 418,
  419, 407,
  420, 419,
  420, 408,
  553, 420,
  421, 409,
  422, 421,
  422, 410,
  423, 422,
  423, 411,
  424, 423,
  424, 412,
  425, 424,
  425, 413,
  426, 425,
  426, 414,
  427, 426,
  427, 415,
  428, 427,
  428, 416,
  429, 428,
  429, 417,
  430, 429,
  430, 418,
  431, 430,
  431, 419,
  432, 431,
  432, 420,
  565, 432,
  854, 421,
  855, 854,
  855, 422,
  856, 855,
  856, 423,
  857, 856,
  857, 424,
  858, 857,
  858, 425,
  859, 858,
  859, 426,
  860, 859,
  860, 427,
  861, 860,
  861, 428,
  862, 861,
  862, 429,
  863, 862,
  863, 430,
  864, 863,
  864, 431,
  865, 864,
  865, 432,
  866, 865,
  433, 434,
  445, 433,
  446, 445,
  434, 435,
  446, 434,
  447, 446,
  435, 436,
  447, 435,
  448, 447,
  436, 437,
  448, 436,
  449, 448,
  437, 438,
  449, 437,
  450, 449,
  438, 439,
  450, 438,
  451, 450,
  439, 440,
  451, 439,
  452, 451,
  440, 441,
  452, 440,
  453, 452,
  441, 442,
  453, 441,
  454, 453,
  442, 443,
  454, 442,
  455, 454,
  443, 444,
  455, 443,
  456, 455,
  444, 1,
  456, 444,
  13, 456,
  457, 445,
  458, 457,
  458, 446,
  459, 458,
  459, 447,
  460, 459,
  460, 448,
  461, 460,
  461, 449,
  462, 461,
  462, 450,
  463, 462,
  463, 451,
  464, 463,
  464, 452,
  465, 464,
  465, 453,
  466, 465,
  466, 454,
  467, 466,
  467, 455,
  468, 467,
  468, 456,
  25, 468,
  469, 457,
  470, 469,
  470, 458,
  471, 470,
  471, 459,
  472, 471,
  472, 460,
  473, 472,
  473, 461,
  474, 473,
  474, 462,
  475, 474,
  475, 463,
  476, 475,
  476, 464,
  477, 476,
  477, 465,
  478, 477,
  478, 466,
  479, 478,
  479, 467,
  480, 479,
  480, 468,
  37, 480,
  481, 469,
  482, 481,
  482, 470,
  483, 482,
  483, 471,
  484, 483,
  484, 472,
  485, 484,
  485, 473,
  486, 485,
  486, 474,
  487, 486,
  487, 475,
  488, 487,
  488, 476,
  489, 488,
  489, 477,
  490, 489,
  490, 478,
  491, 490,
  491, 479,
  492, 491,
  492, 480,
  49, 492,
  493, 481,
  494, 493,
  494, 482,
  495, 494,
  495, 483,
  496, 495,
  496, 484,
  497, 496,
  497, 485,
  498, 497,
  498, 486,
  499, 498,
  499, 487,
  500, 499,
  500, 488,
  501, 500,
  501, 489,
  502, 501,
  502, 490,
  503, 502,
  503, 491,
  504, 503,
  504, 492,
  61, 504,
  505, 493,
  506, 505,
  506, 494,
  507, 506,
  507, 495,
  508, 507,
  508, 496,
  509, 508,
  509, 497,
  510, 509,
  510, 498,
  511, 510,
  511, 499,
  512, 511,
  512, 500,
  513, 512,
  513, 501,
  514, 513,
  514, 502,
  515, 514,
  515, 503,
  516, 515,
  516, 504,
  73, 516,
  517, 505,
  518, 517,
  518, 506,
  519, 518,
  519, 507,
  520, 519,
  520, 508,
  521, 520,
  521, 509,
  522, 521,
  522, 510,
  523, 522,
  523, 511,
  524, 523,
  524, 512,
  525, 524,
  525, 513,
  526, 525,
  526, 514,
  527, 526,
  527, 515,
  528, 527,
  528, 516,
  85, 528,
  529, 517,
  530, 529,
  530, 518,
  531, 530,
  531, 519,
  532, 531,
  532, 520,
  533, 532,
  533, 521,
  534, 533,
  534, 522,
  535, 534,
  535, 523,
  536, 535,
  536, 524,
  537, 536,
  537, 525,
  538, 537,
  538, 526,
  539, 538,
  539, 527,
  540, 539,
  540, 528,
  97, 540,
  541, 529,
  542, 541,
  542, 530,
  543, 542,
  543, 531,
  544, 543,
  544, 532,
  545, 544,
  545, 533,
  546, 545,
  546, 534,
  547, 546,
  547, 535,
  548, 547,
  548, 536,
  549, 548,
  549, 537,
  550, 549,
  550, 538,
  551, 550,
  551, 539,
  552, 551,
  552, 540,
  109, 552,
  553, 541,
  554, 553,
  554, 542,
  555, 554,
  555, 543,
  556, 555,
  556, 544,
  557, 556,
  557, 545,
  558, 557,
  558, 546,
  559, 558,
  559, 547,
  560, 559,
  560, 548,
  561, 560,
  561, 549,
  562, 561,
  562, 550,
  563, 562,
  563, 551,
  564, 563,
  564, 552,
  121, 564,
  565, 553,
  566, 565,
  566, 554,
  567, 566,
  567, 555,
  568, 567,
  568, 556,
  569, 568,
  569, 557,
  570, 569,
  570, 558,
  571, 570,
  571, 559,
  572, 571,
  572, 560,
  573, 572,
  573, 561,
  574, 573,
  574, 562,
  575, 574,
  575, 563,
  576, 575,
  576, 564,
  133, 576,
  866, 565,
  853, 866,
  853, 566,
  852, 853,
  852, 567,
  851, 852,
  851, 568,
  850, 851,
  850, 569,
  849, 850,
  849, 570,
  848, 849,
  848, 571,
  847, 848,
  847, 572,
  846, 847,
  846, 573,
  845, 846,
  845, 574,
  844, 845,
  844, 575,
  843, 844,
  843, 576,
  842, 843,
  577, 2,
  578, 577,
  579, 578,
  580, 579,
  581, 580,
  582, 581,
  583, 582,
  584, 583,
  585, 584,
  586, 585,
  587, 586,
  300, 587,
  588, 3,
  589, 588,
  590, 589,
  591, 590,
  592, 591,
  593, 592,
  594, 593,
  595, 594,
  596, 595,
  597, 596,
  598, 597,
  299, 598,
  599, 4,
  600, 599,
  601, 600,
  602, 601,
  603, 602,
  604, 603,
  605, 604,
  606, 605,
  607, 606,
  608, 607,
  609, 608,
  298, 609,
  610, 5,
  611, 610,
  612, 611,
  613, 612,
  614, 613,
  615, 614,
  616, 615,
  617, 616,
  618, 617,
  619, 618,
  620, 619,
  297, 620,
  621, 6,
  622, 621,
  623, 622,
  624, 623,
  625, 624,
  626, 625,
  627, 626,
  628, 627,
  629, 628,
  630, 629,
  631, 630,
  296, 631,
  632, 7,
  633, 632,
  634, 633,
  635, 634,
  636, 635,
  637, 636,
  638, 637,
  639, 638,
  640, 639,
  641, 640,
  642, 641,
  295, 642,
  643, 8,
  644, 643,
  645, 644,
  646, 645,
  647, 646,
  648, 647,
  649, 648,
  650, 649,
  651, 650,
  652, 651,
  653, 652,
  294, 653,
  654, 9,
  655, 654,
  656, 655,
  657, 656,
  658, 657,
  659, 658,
  660, 659,
  661, 660,
  662, 661,
  663, 662,
  664, 663,
  293, 664,
  665, 10,
  666, 665,
  667, 666,
  668, 667,
  669, 668,
  670, 669,
  671, 670,
  672, 671,
  673, 672,
  674, 673,
  675, 674,
  292, 675,
  676, 11,
  677, 676,
  678, 677,
  679, 678,
  680, 679,
  681, 680,
  682, 681,
  683, 682,
  684, 683,
  685, 684,
  686, 685,
  291, 686,
  687, 12,
  688, 687,
  689, 688,
  690, 689,
  691, 690,
  692, 691,
  693, 692,
  694, 693,
  695, 694,
  696, 695,
  697, 696,
  290, 697,
  444, 577,
  443, 578,
  442, 579,
  441, 580,
  440, 581,
  439, 582,
  438, 583,
  437, 584,
  436, 585,
  435, 586,
  434, 587,
  577, 588,
  578, 589,
  579, 590,
  580, 591,
  581, 592,
  582, 593,
  583, 594,
  584, 595,
  585, 596,
  586, 597,
  587, 598,
  588, 599,
  589, 600,
  590, 601,
  591, 602,
  592, 603,
  593, 604,
  594, 605,
  595, 606,
  596, 607,
  597, 608,
  598, 609,
  599, 610,
  600, 611,
  601, 612,
  602, 613,
  603, 614,
  604, 615,
  605, 616,
  606, 617,
  607, 618,
  608, 619,
  609, 620,
  610, 621,
  611, 622,
  612, 623,
  613, 624,
  614, 625,
  615, 626,
  616, 627,
  617, 628,
  618, 629,
  619, 630,
  620, 631,
  621, 632,
  622, 633,
  623, 634,
  624, 635,
  625, 636,
  626, 637,
  627, 638,
  628, 639,
  629, 640,
  630, 641,
  631, 642,
  632, 643,
  633, 644,
  634, 645,
  635, 646,
  636, 647,
  637, 648,
  638, 649,
  639, 650,
  640, 651,
  641, 652,
  642, 653,
  643, 654,
  644, 655,
  645, 656,
  646, 657,
  647, 658,
  648, 659,
  649, 660,
  650, 661,
  651, 662,
  652, 663,
  653, 664,
  654, 665,
  655, 666,
  656, 667,
  657, 668,
  658, 669,
  659, 670,
  660, 671,
  661, 672,
  662, 673,
  663, 674,
  664, 675,
  665, 676,
  666, 677,
  667, 678,
  668, 679,
  669, 680,
  670, 681,
  671, 682,
  672, 683,
  673, 684,
  674, 685,
  675, 686,
  676, 687,
  677, 688,
  678, 689,
  679, 690,
  680, 691,
  681, 692,
  682, 693,
  683, 694,
  684, 695,
  685, 696,
  686, 697,
  687, 146,
  688, 147,
  689, 148,
  690, 149,
  691, 150,
  692, 151,
  693, 152,
  694, 153,
  695, 154,
  696, 155,
  697, 156,
  711, 710,
  712, 711,
  713, 712,
  714, 713,
  715, 714,
  716, 715,
  717, 716,
  718, 717,
  719, 718,
  720, 719,
  721, 720,
  855, 721,
  723, 722,
  724, 723,
  725, 724,
  726, 725,
  727, 726,
  728, 727,
  729, 728,
  730, 729,
  731, 730,
  732, 731,
  733, 732,
  856, 733,
  735, 734,
  736, 735,
  737, 736,
  738, 737,
  739, 738,
  740, 739,
  741, 740,
  742, 741,
  743, 742,
  744, 743,
  745, 744,
  857, 745,
  747, 746,
  748, 747,
  749, 748,
  750, 749,
  751, 750,
  752, 751,
  753, 752,
  754, 753,
  755, 754,
  756, 755,
  757, 756,
  858, 757,
  759, 758,
  760, 759,
  761, 760,
  762, 761,
  763, 762,
  764, 763,
  765, 764,
  766, 765,
  767, 766,
  768, 767,
  769, 768,
  859, 769,
  771, 770,
  772, 771,
  773, 772,
  774, 773,
  775, 774,
  776, 775,
  777, 776,
  778, 777,
  779, 778,
  780, 779,
  781, 780,
  860, 781,
  783, 782,
  784, 783,
  785, 784,
  786, 785,
  787, 786,
  788, 787,
  789, 788,
  790, 789,
  791, 790,
  792, 791,
  793, 792,
  861, 793,
  795, 794,
  796, 795,
  797, 796,
  798, 797,
  799, 798,
  800, 799,
  801, 800,
  802, 801,
  803, 802,
  804, 803,
  805, 804,
  862, 805,
  807, 806,
  808, 807,
  809, 808,
  810, 809,
  811, 810,
  812, 811,
  813, 812,
  814, 813,
  815, 814,
  816, 815,
  817, 816,
  863, 817,
  819, 818,
  820, 819,
  821, 820,
  822, 821,
  823, 822,
  824, 823,
  825, 824,
  826, 825,
  827, 826,
  828, 827,
  829, 828,
  864, 829,
  831, 830,
  832, 831,
  833, 832,
  834, 833,
  835, 834,
  836, 835,
  837, 836,
  838, 837,
  839, 838,
  840, 839,
  841, 840,
  865, 841,
  699, 711,
  700, 712,
  701, 713,
  702, 714,
  703, 715,
  704, 716,
  705, 717,
  706, 718,
  707, 719,
  708, 720,
  709, 721,
  711, 723,
  712, 724,
  713, 725,
  714, 726,
  715, 727,
  716, 728,
  717, 729,
  718, 730,
  719, 731,
  720, 732,
  721, 733,
  723, 735,
  724, 736,
  725, 737,
  726, 738,
  727, 739,
  728, 740,
  729, 741,
  730, 742,
  731, 743,
  732, 744,
  733, 745,
  735, 747,
  736, 748,
  737, 749,
  738, 750,
  739, 751,
  740, 752,
  741, 753,
  742, 754,
  743, 755,
  744, 756,
  745, 757,
  747, 759,
  748, 760,
  749, 761,
  750, 762,
  751, 763,
  752, 764,
  753, 765,
  754, 766,
  755, 767,
  756, 768,
  757, 769,
  759, 771,
  760, 772,
  761, 773,
  762, 774,
  763, 775,
  764, 776,
  765, 777,
  766, 778,
  767, 779,
  768, 780,
  769, 781,
  771, 783,
  772, 784,
  773, 785,
  774, 786,
  775, 787,
  776, 788,
  777, 789,
  778, 790,
  779, 791,
  780, 792,
  781, 793,
  783, 795,
  784, 796,
  785, 797,
  786, 798,
  787, 799,
  788, 800,
  789, 801,
  790, 802,
  791, 803,
  792, 804,
  793, 805,
  795, 807,
  796, 808,
  797, 809,
  798, 810,
  799, 811,
  800, 812,
  801, 813,
  802, 814,
  803, 815,
  804, 816,
  805, 817,
  807, 819,
  808, 820,
  809, 821,
  810, 822,
  811, 823,
  812, 824,
  813, 825,
  814, 826,
  815, 827,
  816, 828,
  817, 829,
  819, 831,
  820, 832,
  821, 833,
  822, 834,
  823, 835,
  824, 836,
  825, 837,
  826, 838,
  827, 839,
  828, 840,
  829, 841,
  831, 843,
  832, 844,
  833, 845,
  834, 846,
  835, 847,
  836, 848,
  837, 849,
  838, 850,
  839, 851,
  840, 852,
  841, 853 ;

 dynamics_face_edges =
  2, 3, 5, 1,
  5, 6, 8, 4,
  8, 9, 11, 7,
  11, 12, 14, 10,
  14, 15, 17, 13,
  17, 18, 20, 16,
  20, 21, 23, 19,
  23, 24, 26, 22,
  26, 27, 29, 25,
  29, 30, 32, 28,
  32, 33, 35, 31,
  35, 36, 302, 34,
  37, 38, 39, 3,
  39, 40, 41, 6,
  41, 42, 43, 9,
  43, 44, 45, 12,
  45, 46, 47, 15,
  47, 48, 49, 18,
  49, 50, 51, 21,
  51, 52, 53, 24,
  53, 54, 55, 27,
  55, 56, 57, 30,
  57, 58, 59, 33,
  59, 60, 337, 36,
  61, 62, 63, 38,
  63, 64, 65, 40,
  65, 66, 67, 42,
  67, 68, 69, 44,
  69, 70, 71, 46,
  71, 72, 73, 48,
  73, 74, 75, 50,
  75, 76, 77, 52,
  77, 78, 79, 54,
  79, 80, 81, 56,
  81, 82, 83, 58,
  83, 84, 361, 60,
  85, 86, 87, 62,
  87, 88, 89, 64,
  89, 90, 91, 66,
  91, 92, 93, 68,
  93, 94, 95, 70,
  95, 96, 97, 72,
  97, 98, 99, 74,
  99, 100, 101, 76,
  101, 102, 103, 78,
  103, 104, 105, 80,
  105, 106, 107, 82,
  107, 108, 385, 84,
  109, 110, 111, 86,
  111, 112, 113, 88,
  113, 114, 115, 90,
  115, 116, 117, 92,
  117, 118, 119, 94,
  119, 120, 121, 96,
  121, 122, 123, 98,
  123, 124, 125, 100,
  125, 126, 127, 102,
  127, 128, 129, 104,
  129, 130, 131, 106,
  131, 132, 409, 108,
  133, 134, 135, 110,
  135, 136, 137, 112,
  137, 138, 139, 114,
  139, 140, 141, 116,
  141, 142, 143, 118,
  143, 144, 145, 120,
  145, 146, 147, 122,
  147, 148, 149, 124,
  149, 150, 151, 126,
  151, 152, 153, 128,
  153, 154, 155, 130,
  155, 156, 433, 132,
  157, 158, 159, 134,
  159, 160, 161, 136,
  161, 162, 163, 138,
  163, 164, 165, 140,
  165, 166, 167, 142,
  167, 168, 169, 144,
  169, 170, 171, 146,
  171, 172, 173, 148,
  173, 174, 175, 150,
  175, 176, 177, 152,
  177, 178, 179, 154,
  179, 180, 457, 156,
  181, 182, 183, 158,
  183, 184, 185, 160,
  185, 186, 187, 162,
  187, 188, 189, 164,
  189, 190, 191, 166,
  191, 192, 193, 168,
  193, 194, 195, 170,
  195, 196, 197, 172,
  197, 198, 199, 174,
  199, 200, 201, 176,
  201, 202, 203, 178,
  203, 204, 481, 180,
  205, 206, 207, 182,
  207, 208, 209, 184,
  209, 210, 211, 186,
  211, 212, 213, 188,
  213, 214, 215, 190,
  215, 216, 217, 192,
  217, 218, 219, 194,
  219, 220, 221, 196,
  221, 222, 223, 198,
  223, 224, 225, 200,
  225, 226, 227, 202,
  227, 228, 505, 204,
  229, 230, 231, 206,
  231, 232, 233, 208,
  233, 234, 235, 210,
  235, 236, 237, 212,
  237, 238, 239, 214,
  239, 240, 241, 216,
  241, 242, 243, 218,
  243, 244, 245, 220,
  245, 246, 247, 222,
  247, 248, 249, 224,
  249, 250, 251, 226,
  251, 252, 529, 228,
  253, 254, 255, 230,
  255, 256, 257, 232,
  257, 258, 259, 234,
  259, 260, 261, 236,
  261, 262, 263, 238,
  263, 264, 265, 240,
  265, 266, 267, 242,
  267, 268, 269, 244,
  269, 270, 271, 246,
  271, 272, 273, 248,
  273, 274, 275, 250,
  275, 276, 553, 252,
  277, 278, 279, 254,
  279, 280, 281, 256,
  281, 282, 283, 258,
  283, 284, 285, 260,
  285, 286, 287, 262,
  287, 288, 289, 264,
  289, 290, 291, 266,
  291, 292, 293, 268,
  293, 294, 295, 270,
  295, 296, 297, 272,
  297, 298, 299, 274,
  299, 300, 577, 276,
  302, 303, 305, 301,
  305, 306, 308, 304,
  308, 309, 311, 307,
  311, 312, 314, 310,
  314, 315, 317, 313,
  317, 318, 320, 316,
  320, 321, 323, 319,
  323, 324, 326, 322,
  326, 327, 329, 325,
  329, 330, 332, 328,
  332, 333, 335, 331,
  335, 336, 602, 334,
  337, 338, 339, 303,
  339, 340, 341, 306,
  341, 342, 343, 309,
  343, 344, 345, 312,
  345, 346, 347, 315,
  347, 348, 349, 318,
  349, 350, 351, 321,
  351, 352, 353, 324,
  353, 354, 355, 327,
  355, 356, 357, 330,
  357, 358, 359, 333,
  359, 360, 637, 336,
  361, 362, 363, 338,
  363, 364, 365, 340,
  365, 366, 367, 342,
  367, 368, 369, 344,
  369, 370, 371, 346,
  371, 372, 373, 348,
  373, 374, 375, 350,
  375, 376, 377, 352,
  377, 378, 379, 354,
  379, 380, 381, 356,
  381, 382, 383, 358,
  383, 384, 661, 360,
  385, 386, 387, 362,
  387, 388, 389, 364,
  389, 390, 391, 366,
  391, 392, 393, 368,
  393, 394, 395, 370,
  395, 396, 397, 372,
  397, 398, 399, 374,
  399, 400, 401, 376,
  401, 402, 403, 378,
  403, 404, 405, 380,
  405, 406, 407, 382,
  407, 408, 685, 384,
  409, 410, 411, 386,
  411, 412, 413, 388,
  413, 414, 415, 390,
  415, 416, 417, 392,
  417, 418, 419, 394,
  419, 420, 421, 396,
  421, 422, 423, 398,
  423, 424, 425, 400,
  425, 426, 427, 402,
  427, 428, 429, 404,
  429, 430, 431, 406,
  431, 432, 709, 408,
  433, 434, 435, 410,
  435, 436, 437, 412,
  437, 438, 439, 414,
  439, 440, 441, 416,
  441, 442, 443, 418,
  443, 444, 445, 420,
  445, 446, 447, 422,
  447, 448, 449, 424,
  449, 450, 451, 426,
  451, 452, 453, 428,
  453, 454, 455, 430,
  455, 456, 733, 432,
  457, 458, 459, 434,
  459, 460, 461, 436,
  461, 462, 463, 438,
  463, 464, 465, 440,
  465, 466, 467, 442,
  467, 468, 469, 444,
  469, 470, 471, 446,
  471, 472, 473, 448,
  473, 474, 475, 450,
  475, 476, 477, 452,
  477, 478, 479, 454,
  479, 480, 757, 456,
  481, 482, 483, 458,
  483, 484, 485, 460,
  485, 486, 487, 462,
  487, 488, 489, 464,
  489, 490, 491, 466,
  491, 492, 493, 468,
  493, 494, 495, 470,
  495, 496, 497, 472,
  497, 498, 499, 474,
  499, 500, 501, 476,
  501, 502, 503, 478,
  503, 504, 781, 480,
  505, 506, 507, 482,
  507, 508, 509, 484,
  509, 510, 511, 486,
  511, 512, 513, 488,
  513, 514, 515, 490,
  515, 516, 517, 492,
  517, 518, 519, 494,
  519, 520, 521, 496,
  521, 522, 523, 498,
  523, 524, 525, 500,
  525, 526, 527, 502,
  527, 528, 805, 504,
  529, 530, 531, 506,
  531, 532, 533, 508,
  533, 534, 535, 510,
  535, 536, 537, 512,
  537, 538, 539, 514,
  539, 540, 541, 516,
  541, 542, 543, 518,
  543, 544, 545, 520,
  545, 546, 547, 522,
  547, 548, 549, 524,
  549, 550, 551, 526,
  551, 552, 829, 528,
  553, 554, 555, 530,
  555, 556, 557, 532,
  557, 558, 559, 534,
  559, 560, 561, 536,
  561, 562, 563, 538,
  563, 564, 565, 540,
  565, 566, 567, 542,
  567, 568, 569, 544,
  569, 570, 571, 546,
  571, 572, 573, 548,
  573, 574, 575, 550,
  575, 576, 853, 552,
  577, 578, 579, 554,
  579, 580, 581, 556,
  581, 582, 583, 558,
  583, 584, 585, 560,
  585, 586, 587, 562,
  587, 588, 589, 564,
  589, 590, 591, 566,
  591, 592, 593, 568,
  593, 594, 595, 570,
  595, 596, 597, 572,
  597, 598, 599, 574,
  599, 600, 877, 576,
  603, 605, 601, 602,
  606, 608, 604, 605,
  609, 611, 607, 608,
  612, 614, 610, 611,
  615, 617, 613, 614,
  618, 620, 616, 617,
  621, 623, 619, 620,
  624, 626, 622, 623,
  627, 629, 625, 626,
  630, 632, 628, 629,
  633, 635, 631, 632,
  636, 902, 634, 635,
  638, 639, 603, 637,
  640, 641, 606, 639,
  642, 643, 609, 641,
  644, 645, 612, 643,
  646, 647, 615, 645,
  648, 649, 618, 647,
  650, 651, 621, 649,
  652, 653, 624, 651,
  654, 655, 627, 653,
  656, 657, 630, 655,
  658, 659, 633, 657,
  660, 937, 636, 659,
  662, 663, 638, 661,
  664, 665, 640, 663,
  666, 667, 642, 665,
  668, 669, 644, 667,
  670, 671, 646, 669,
  672, 673, 648, 671,
  674, 675, 650, 673,
  676, 677, 652, 675,
  678, 679, 654, 677,
  680, 681, 656, 679,
  682, 683, 658, 681,
  684, 961, 660, 683,
  686, 687, 662, 685,
  688, 689, 664, 687,
  690, 691, 666, 689,
  692, 693, 668, 691,
  694, 695, 670, 693,
  696, 697, 672, 695,
  698, 699, 674, 697,
  700, 701, 676, 699,
  702, 703, 678, 701,
  704, 705, 680, 703,
  706, 707, 682, 705,
  708, 985, 684, 707,
  710, 711, 686, 709,
  712, 713, 688, 711,
  714, 715, 690, 713,
  716, 717, 692, 715,
  718, 719, 694, 717,
  720, 721, 696, 719,
  722, 723, 698, 721,
  724, 725, 700, 723,
  726, 727, 702, 725,
  728, 729, 704, 727,
  730, 731, 706, 729,
  732, 1009, 708, 731,
  734, 735, 710, 733,
  736, 737, 712, 735,
  738, 739, 714, 737,
  740, 741, 716, 739,
  742, 743, 718, 741,
  744, 745, 720, 743,
  746, 747, 722, 745,
  748, 749, 724, 747,
  750, 751, 726, 749,
  752, 753, 728, 751,
  754, 755, 730, 753,
  756, 1033, 732, 755,
  758, 759, 734, 757,
  760, 761, 736, 759,
  762, 763, 738, 761,
  764, 765, 740, 763,
  766, 767, 742, 765,
  768, 769, 744, 767,
  770, 771, 746, 769,
  772, 773, 748, 771,
  774, 775, 750, 773,
  776, 777, 752, 775,
  778, 779, 754, 777,
  780, 1057, 756, 779,
  782, 783, 758, 781,
  784, 785, 760, 783,
  786, 787, 762, 785,
  788, 789, 764, 787,
  790, 791, 766, 789,
  792, 793, 768, 791,
  794, 795, 770, 793,
  796, 797, 772, 795,
  798, 799, 774, 797,
  800, 801, 776, 799,
  802, 803, 778, 801,
  804, 1081, 780, 803,
  806, 807, 782, 805,
  808, 809, 784, 807,
  810, 811, 786, 809,
  812, 813, 788, 811,
  814, 815, 790, 813,
  816, 817, 792, 815,
  818, 819, 794, 817,
  820, 821, 796, 819,
  822, 823, 798, 821,
  824, 825, 800, 823,
  826, 827, 802, 825,
  828, 1105, 804, 827,
  830, 831, 806, 829,
  832, 833, 808, 831,
  834, 835, 810, 833,
  836, 837, 812, 835,
  838, 839, 814, 837,
  840, 841, 816, 839,
  842, 843, 818, 841,
  844, 845, 820, 843,
  846, 847, 822, 845,
  848, 849, 824, 847,
  850, 851, 826, 849,
  852, 1129, 828, 851,
  854, 855, 830, 853,
  856, 857, 832, 855,
  858, 859, 834, 857,
  860, 861, 836, 859,
  862, 863, 838, 861,
  864, 865, 840, 863,
  866, 867, 842, 865,
  868, 869, 844, 867,
  870, 871, 846, 869,
  872, 873, 848, 871,
  874, 875, 850, 873,
  876, 1153, 852, 875,
  878, 879, 854, 877,
  880, 881, 856, 879,
  882, 883, 858, 881,
  884, 885, 860, 883,
  886, 887, 862, 885,
  888, 889, 864, 887,
  890, 891, 866, 889,
  892, 893, 868, 891,
  894, 895, 870, 893,
  896, 897, 872, 895,
  898, 899, 874, 897,
  900, 1177, 876, 899,
  903, 905, 901, 902,
  906, 908, 904, 905,
  909, 911, 907, 908,
  912, 914, 910, 911,
  915, 917, 913, 914,
  918, 920, 916, 917,
  921, 923, 919, 920,
  924, 926, 922, 923,
  927, 929, 925, 926,
  930, 932, 928, 929,
  933, 935, 931, 932,
  936, 2, 934, 935,
  938, 939, 903, 937,
  940, 941, 906, 939,
  942, 943, 909, 941,
  944, 945, 912, 943,
  946, 947, 915, 945,
  948, 949, 918, 947,
  950, 951, 921, 949,
  952, 953, 924, 951,
  954, 955, 927, 953,
  956, 957, 930, 955,
  958, 959, 933, 957,
  960, 37, 936, 959,
  962, 963, 938, 961,
  964, 965, 940, 963,
  966, 967, 942, 965,
  968, 969, 944, 967,
  970, 971, 946, 969,
  972, 973, 948, 971,
  974, 975, 950, 973,
  976, 977, 952, 975,
  978, 979, 954, 977,
  980, 981, 956, 979,
  982, 983, 958, 981,
  984, 61, 960, 983,
  986, 987, 962, 985,
  988, 989, 964, 987,
  990, 991, 966, 989,
  992, 993, 968, 991,
  994, 995, 970, 993,
  996, 997, 972, 995,
  998, 999, 974, 997,
  1000, 1001, 976, 999,
  1002, 1003, 978, 1001,
  1004, 1005, 980, 1003,
  1006, 1007, 982, 1005,
  1008, 85, 984, 1007,
  1010, 1011, 986, 1009,
  1012, 1013, 988, 1011,
  1014, 1015, 990, 1013,
  1016, 1017, 992, 1015,
  1018, 1019, 994, 1017,
  1020, 1021, 996, 1019,
  1022, 1023, 998, 1021,
  1024, 1025, 1000, 1023,
  1026, 1027, 1002, 1025,
  1028, 1029, 1004, 1027,
  1030, 1031, 1006, 1029,
  1032, 109, 1008, 1031,
  1034, 1035, 1010, 1033,
  1036, 1037, 1012, 1035,
  1038, 1039, 1014, 1037,
  1040, 1041, 1016, 1039,
  1042, 1043, 1018, 1041,
  1044, 1045, 1020, 1043,
  1046, 1047, 1022, 1045,
  1048, 1049, 1024, 1047,
  1050, 1051, 1026, 1049,
  1052, 1053, 1028, 1051,
  1054, 1055, 1030, 1053,
  1056, 133, 1032, 1055,
  1058, 1059, 1034, 1057,
  1060, 1061, 1036, 1059,
  1062, 1063, 1038, 1061,
  1064, 1065, 1040, 1063,
  1066, 1067, 1042, 1065,
  1068, 1069, 1044, 1067,
  1070, 1071, 1046, 1069,
  1072, 1073, 1048, 1071,
  1074, 1075, 1050, 1073,
  1076, 1077, 1052, 1075,
  1078, 1079, 1054, 1077,
  1080, 157, 1056, 1079,
  1082, 1083, 1058, 1081,
  1084, 1085, 1060, 1083,
  1086, 1087, 1062, 1085,
  1088, 1089, 1064, 1087,
  1090, 1091, 1066, 1089,
  1092, 1093, 1068, 1091,
  1094, 1095, 1070, 1093,
  1096, 1097, 1072, 1095,
  1098, 1099, 1074, 1097,
  1100, 1101, 1076, 1099,
  1102, 1103, 1078, 1101,
  1104, 181, 1080, 1103,
  1106, 1107, 1082, 1105,
  1108, 1109, 1084, 1107,
  1110, 1111, 1086, 1109,
  1112, 1113, 1088, 1111,
  1114, 1115, 1090, 1113,
  1116, 1117, 1092, 1115,
  1118, 1119, 1094, 1117,
  1120, 1121, 1096, 1119,
  1122, 1123, 1098, 1121,
  1124, 1125, 1100, 1123,
  1126, 1127, 1102, 1125,
  1128, 205, 1104, 1127,
  1130, 1131, 1106, 1129,
  1132, 1133, 1108, 1131,
  1134, 1135, 1110, 1133,
  1136, 1137, 1112, 1135,
  1138, 1139, 1114, 1137,
  1140, 1141, 1116, 1139,
  1142, 1143, 1118, 1141,
  1144, 1145, 1120, 1143,
  1146, 1147, 1122, 1145,
  1148, 1149, 1124, 1147,
  1150, 1151, 1126, 1149,
  1152, 229, 1128, 1151,
  1154, 1155, 1130, 1153,
  1156, 1157, 1132, 1155,
  1158, 1159, 1134, 1157,
  1160, 1161, 1136, 1159,
  1162, 1163, 1138, 1161,
  1164, 1165, 1140, 1163,
  1166, 1167, 1142, 1165,
  1168, 1169, 1144, 1167,
  1170, 1171, 1146, 1169,
  1172, 1173, 1148, 1171,
  1174, 1175, 1150, 1173,
  1176, 253, 1152, 1175,
  1178, 1179, 1154, 1177,
  1180, 1181, 1156, 1179,
  1182, 1183, 1158, 1181,
  1184, 1185, 1160, 1183,
  1186, 1187, 1162, 1185,
  1188, 1189, 1164, 1187,
  1190, 1191, 1166, 1189,
  1192, 1193, 1168, 1191,
  1194, 1195, 1170, 1193,
  1196, 1197, 1172, 1195,
  1198, 1199, 1174, 1197,
  1200, 277, 1176, 1199,
  934, 1, 1201, 1333,
  931, 1333, 1202, 1334,
  928, 1334, 1203, 1335,
  925, 1335, 1204, 1336,
  922, 1336, 1205, 1337,
  919, 1337, 1206, 1338,
  916, 1338, 1207, 1339,
  913, 1339, 1208, 1340,
  910, 1340, 1209, 1341,
  907, 1341, 1210, 1342,
  904, 1342, 1211, 1343,
  901, 1343, 1212, 634,
  1201, 4, 1213, 1344,
  1202, 1344, 1214, 1345,
  1203, 1345, 1215, 1346,
  1204, 1346, 1216, 1347,
  1205, 1347, 1217, 1348,
  1206, 1348, 1218, 1349,
  1207, 1349, 1219, 1350,
  1208, 1350, 1220, 1351,
  1209, 1351, 1221, 1352,
  1210, 1352, 1222, 1353,
  1211, 1353, 1223, 1354,
  1212, 1354, 1224, 631,
  1213, 7, 1225, 1355,
  1214, 1355, 1226, 1356,
  1215, 1356, 1227, 1357,
  1216, 1357, 1228, 1358,
  1217, 1358, 1229, 1359,
  1218, 1359, 1230, 1360,
  1219, 1360, 1231, 1361,
  1220, 1361, 1232, 1362,
  1221, 1362, 1233, 1363,
  1222, 1363, 1234, 1364,
  1223, 1364, 1235, 1365,
  1224, 1365, 1236, 628,
  1225, 10, 1237, 1366,
  1226, 1366, 1238, 1367,
  1227, 1367, 1239, 1368,
  1228, 1368, 1240, 1369,
  1229, 1369, 1241, 1370,
  1230, 1370, 1242, 1371,
  1231, 1371, 1243, 1372,
  1232, 1372, 1244, 1373,
  1233, 1373, 1245, 1374,
  1234, 1374, 1246, 1375,
  1235, 1375, 1247, 1376,
  1236, 1376, 1248, 625,
  1237, 13, 1249, 1377,
  1238, 1377, 1250, 1378,
  1239, 1378, 1251, 1379,
  1240, 1379, 1252, 1380,
  1241, 1380, 1253, 1381,
  1242, 1381, 1254, 1382,
  1243, 1382, 1255, 1383,
  1244, 1383, 1256, 1384,
  1245, 1384, 1257, 1385,
  1246, 1385, 1258, 1386,
  1247, 1386, 1259, 1387,
  1248, 1387, 1260, 622,
  1249, 16, 1261, 1388,
  1250, 1388, 1262, 1389,
  1251, 1389, 1263, 1390,
  1252, 1390, 1264, 1391,
  1253, 1391, 1265, 1392,
  1254, 1392, 1266, 1393,
  1255, 1393, 1267, 1394,
  1256, 1394, 1268, 1395,
  1257, 1395, 1269, 1396,
  1258, 1396, 1270, 1397,
  1259, 1397, 1271, 1398,
  1260, 1398, 1272, 619,
  1261, 19, 1273, 1399,
  1262, 1399, 1274, 1400,
  1263, 1400, 1275, 1401,
  1264, 1401, 1276, 1402,
  1265, 1402, 1277, 1403,
  1266, 1403, 1278, 1404,
  1267, 1404, 1279, 1405,
  1268, 1405, 1280, 1406,
  1269, 1406, 1281, 1407,
  1270, 1407, 1282, 1408,
  1271, 1408, 1283, 1409,
  1272, 1409, 1284, 616,
  1273, 22, 1285, 1410,
  1274, 1410, 1286, 1411,
  1275, 1411, 1287, 1412,
  1276, 1412, 1288, 1413,
  1277, 1413, 1289, 1414,
  1278, 1414, 1290, 1415,
  1279, 1415, 1291, 1416,
  1280, 1416, 1292, 1417,
  1281, 1417, 1293, 1418,
  1282, 1418, 1294, 1419,
  1283, 1419, 1295, 1420,
  1284, 1420, 1296, 613,
  1285, 25, 1297, 1421,
  1286, 1421, 1298, 1422,
  1287, 1422, 1299, 1423,
  1288, 1423, 1300, 1424,
  1289, 1424, 1301, 1425,
  1290, 1425, 1302, 1426,
  1291, 1426, 1303, 1427,
  1292, 1427, 1304, 1428,
  1293, 1428, 1305, 1429,
  1294, 1429, 1306, 1430,
  1295, 1430, 1307, 1431,
  1296, 1431, 1308, 610,
  1297, 28, 1309, 1432,
  1298, 1432, 1310, 1433,
  1299, 1433, 1311, 1434,
  1300, 1434, 1312, 1435,
  1301, 1435, 1313, 1436,
  1302, 1436, 1314, 1437,
  1303, 1437, 1315, 1438,
  1304, 1438, 1316, 1439,
  1305, 1439, 1317, 1440,
  1306, 1440, 1318, 1441,
  1307, 1441, 1319, 1442,
  1308, 1442, 1320, 607,
  1309, 31, 1321, 1443,
  1310, 1443, 1322, 1444,
  1311, 1444, 1323, 1445,
  1312, 1445, 1324, 1446,
  1313, 1446, 1325, 1447,
  1314, 1447, 1326, 1448,
  1315, 1448, 1327, 1449,
  1316, 1449, 1328, 1450,
  1317, 1450, 1329, 1451,
  1318, 1451, 1330, 1452,
  1319, 1452, 1331, 1453,
  1320, 1453, 1332, 604,
  1321, 34, 301, 1454,
  1322, 1454, 304, 1455,
  1323, 1455, 307, 1456,
  1324, 1456, 310, 1457,
  1325, 1457, 313, 1458,
  1326, 1458, 316, 1459,
  1327, 1459, 319, 1460,
  1328, 1460, 322, 1461,
  1329, 1461, 325, 1462,
  1330, 1462, 328, 1463,
  1331, 1463, 331, 1464,
  1332, 1464, 334, 601,
  300, 1465, 1597, 578,
  1597, 1466, 1598, 580,
  1598, 1467, 1599, 582,
  1599, 1468, 1600, 584,
  1600, 1469, 1601, 586,
  1601, 1470, 1602, 588,
  1602, 1471, 1603, 590,
  1603, 1472, 1604, 592,
  1604, 1473, 1605, 594,
  1605, 1474, 1606, 596,
  1606, 1475, 1607, 598,
  1607, 1476, 878, 600,
  298, 1477, 1608, 1465,
  1608, 1478, 1609, 1466,
  1609, 1479, 1610, 1467,
  1610, 1480, 1611, 1468,
  1611, 1481, 1612, 1469,
  1612, 1482, 1613, 1470,
  1613, 1483, 1614, 1471,
  1614, 1484, 1615, 1472,
  1615, 1485, 1616, 1473,
  1616, 1486, 1617, 1474,
  1617, 1487, 1618, 1475,
  1618, 1488, 880, 1476,
  296, 1489, 1619, 1477,
  1619, 1490, 1620, 1478,
  1620, 1491, 1621, 1479,
  1621, 1492, 1622, 1480,
  1622, 1493, 1623, 1481,
  1623, 1494, 1624, 1482,
  1624, 1495, 1625, 1483,
  1625, 1496, 1626, 1484,
  1626, 1497, 1627, 1485,
  1627, 1498, 1628, 1486,
  1628, 1499, 1629, 1487,
  1629, 1500, 882, 1488,
  294, 1501, 1630, 1489,
  1630, 1502, 1631, 1490,
  1631, 1503, 1632, 1491,
  1632, 1504, 1633, 1492,
  1633, 1505, 1634, 1493,
  1634, 1506, 1635, 1494,
  1635, 1507, 1636, 1495,
  1636, 1508, 1637, 1496,
  1637, 1509, 1638, 1497,
  1638, 1510, 1639, 1498,
  1639, 1511, 1640, 1499,
  1640, 1512, 884, 1500,
  292, 1513, 1641, 1501,
  1641, 1514, 1642, 1502,
  1642, 1515, 1643, 1503,
  1643, 1516, 1644, 1504,
  1644, 1517, 1645, 1505,
  1645, 1518, 1646, 1506,
  1646, 1519, 1647, 1507,
  1647, 1520, 1648, 1508,
  1648, 1521, 1649, 1509,
  1649, 1522, 1650, 1510,
  1650, 1523, 1651, 1511,
  1651, 1524, 886, 1512,
  290, 1525, 1652, 1513,
  1652, 1526, 1653, 1514,
  1653, 1527, 1654, 1515,
  1654, 1528, 1655, 1516,
  1655, 1529, 1656, 1517,
  1656, 1530, 1657, 1518,
  1657, 1531, 1658, 1519,
  1658, 1532, 1659, 1520,
  1659, 1533, 1660, 1521,
  1660, 1534, 1661, 1522,
  1661, 1535, 1662, 1523,
  1662, 1536, 888, 1524,
  288, 1537, 1663, 1525,
  1663, 1538, 1664, 1526,
  1664, 1539, 1665, 1527,
  1665, 1540, 1666, 1528,
  1666, 1541, 1667, 1529,
  1667, 1542, 1668, 1530,
  1668, 1543, 1669, 1531,
  1669, 1544, 1670, 1532,
  1670, 1545, 1671, 1533,
  1671, 1546, 1672, 1534,
  1672, 1547, 1673, 1535,
  1673, 1548, 890, 1536,
  286, 1549, 1674, 1537,
  1674, 1550, 1675, 1538,
  1675, 1551, 1676, 1539,
  1676, 1552, 1677, 1540,
  1677, 1553, 1678, 1541,
  1678, 1554, 1679, 1542,
  1679, 1555, 1680, 1543,
  1680, 1556, 1681, 1544,
  1681, 1557, 1682, 1545,
  1682, 1558, 1683, 1546,
  1683, 1559, 1684, 1547,
  1684, 1560, 892, 1548,
  284, 1561, 1685, 1549,
  1685, 1562, 1686, 1550,
  1686, 1563, 1687, 1551,
  1687, 1564, 1688, 1552,
  1688, 1565, 1689, 1553,
  1689, 1566, 1690, 1554,
  1690, 1567, 1691, 1555,
  1691, 1568, 1692, 1556,
  1692, 1569, 1693, 1557,
  1693, 1570, 1694, 1558,
  1694, 1571, 1695, 1559,
  1695, 1572, 894, 1560,
  282, 1573, 1696, 1561,
  1696, 1574, 1697, 1562,
  1697, 1575, 1698, 1563,
  1698, 1576, 1699, 1564,
  1699, 1577, 1700, 1565,
  1700, 1578, 1701, 1566,
  1701, 1579, 1702, 1567,
  1702, 1580, 1703, 1568,
  1703, 1581, 1704, 1569,
  1704, 1582, 1705, 1570,
  1705, 1583, 1706, 1571,
  1706, 1584, 896, 1572,
  280, 1585, 1707, 1573,
  1707, 1586, 1708, 1574,
  1708, 1587, 1709, 1575,
  1709, 1588, 1710, 1576,
  1710, 1589, 1711, 1577,
  1711, 1590, 1712, 1578,
  1712, 1591, 1713, 1579,
  1713, 1592, 1714, 1580,
  1714, 1593, 1715, 1581,
  1715, 1594, 1716, 1582,
  1716, 1595, 1717, 1583,
  1717, 1596, 898, 1584,
  278, 1200, 1718, 1585,
  1718, 1198, 1719, 1586,
  1719, 1196, 1720, 1587,
  1720, 1194, 1721, 1588,
  1721, 1192, 1722, 1589,
  1722, 1190, 1723, 1590,
  1723, 1188, 1724, 1591,
  1724, 1186, 1725, 1592,
  1725, 1184, 1726, 1593,
  1726, 1182, 1727, 1594,
  1727, 1180, 1728, 1595,
  1728, 1178, 900, 1596 ;

 dynamics_face_links =
  444, 13, 2, 577,
  1, 14, 3, 589,
  2, 15, 4, 601,
  3, 16, 5, 613,
  4, 17, 6, 625,
  5, 18, 7, 637,
  6, 19, 8, 649,
  7, 20, 9, 661,
  8, 21, 10, 673,
  9, 22, 11, 685,
  10, 23, 12, 697,
  11, 24, 145, 709,
  456, 25, 14, 1,
  13, 26, 15, 2,
  14, 27, 16, 3,
  15, 28, 17, 4,
  16, 29, 18, 5,
  17, 30, 19, 6,
  18, 31, 20, 7,
  19, 32, 21, 8,
  20, 33, 22, 9,
  21, 34, 23, 10,
  22, 35, 24, 11,
  23, 36, 157, 12,
  468, 37, 26, 13,
  25, 38, 27, 14,
  26, 39, 28, 15,
  27, 40, 29, 16,
  28, 41, 30, 17,
  29, 42, 31, 18,
  30, 43, 32, 19,
  31, 44, 33, 20,
  32, 45, 34, 21,
  33, 46, 35, 22,
  34, 47, 36, 23,
  35, 48, 169, 24,
  480, 49, 38, 25,
  37, 50, 39, 26,
  38, 51, 40, 27,
  39, 52, 41, 28,
  40, 53, 42, 29,
  41, 54, 43, 30,
  42, 55, 44, 31,
  43, 56, 45, 32,
  44, 57, 46, 33,
  45, 58, 47, 34,
  46, 59, 48, 35,
  47, 60, 181, 36,
  492, 61, 50, 37,
  49, 62, 51, 38,
  50, 63, 52, 39,
  51, 64, 53, 40,
  52, 65, 54, 41,
  53, 66, 55, 42,
  54, 67, 56, 43,
  55, 68, 57, 44,
  56, 69, 58, 45,
  57, 70, 59, 46,
  58, 71, 60, 47,
  59, 72, 193, 48,
  504, 73, 62, 49,
  61, 74, 63, 50,
  62, 75, 64, 51,
  63, 76, 65, 52,
  64, 77, 66, 53,
  65, 78, 67, 54,
  66, 79, 68, 55,
  67, 80, 69, 56,
  68, 81, 70, 57,
  69, 82, 71, 58,
  70, 83, 72, 59,
  71, 84, 205, 60,
  516, 85, 74, 61,
  73, 86, 75, 62,
  74, 87, 76, 63,
  75, 88, 77, 64,
  76, 89, 78, 65,
  77, 90, 79, 66,
  78, 91, 80, 67,
  79, 92, 81, 68,
  80, 93, 82, 69,
  81, 94, 83, 70,
  82, 95, 84, 71,
  83, 96, 217, 72,
  528, 97, 86, 73,
  85, 98, 87, 74,
  86, 99, 88, 75,
  87, 100, 89, 76,
  88, 101, 90, 77,
  89, 102, 91, 78,
  90, 103, 92, 79,
  91, 104, 93, 80,
  92, 105, 94, 81,
  93, 106, 95, 82,
  94, 107, 96, 83,
  95, 108, 229, 84,
  540, 109, 98, 85,
  97, 110, 99, 86,
  98, 111, 100, 87,
  99, 112, 101, 88,
  100, 113, 102, 89,
  101, 114, 103, 90,
  102, 115, 104, 91,
  103, 116, 105, 92,
  104, 117, 106, 93,
  105, 118, 107, 94,
  106, 119, 108, 95,
  107, 120, 241, 96,
  552, 121, 110, 97,
  109, 122, 111, 98,
  110, 123, 112, 99,
  111, 124, 113, 100,
  112, 125, 114, 101,
  113, 126, 115, 102,
  114, 127, 116, 103,
  115, 128, 117, 104,
  116, 129, 118, 105,
  117, 130, 119, 106,
  118, 131, 120, 107,
  119, 132, 253, 108,
  564, 133, 122, 109,
  121, 134, 123, 110,
  122, 135, 124, 111,
  123, 136, 125, 112,
  124, 137, 126, 113,
  125, 138, 127, 114,
  126, 139, 128, 115,
  127, 140, 129, 116,
  128, 141, 130, 117,
  129, 142, 131, 118,
  130, 143, 132, 119,
  131, 144, 265, 120,
  576, 853, 134, 121,
  133, 841, 135, 122,
  134, 829, 136, 123,
  135, 817, 137, 124,
  136, 805, 138, 125,
  137, 793, 139, 126,
  138, 781, 140, 127,
  139, 769, 141, 128,
  140, 757, 142, 129,
  141, 745, 143, 130,
  142, 733, 144, 131,
  143, 721, 277, 132,
  12, 157, 146, 709,
  145, 158, 147, 710,
  146, 159, 148, 711,
  147, 160, 149, 712,
  148, 161, 150, 713,
  149, 162, 151, 714,
  150, 163, 152, 715,
  151, 164, 153, 716,
  152, 165, 154, 717,
  153, 166, 155, 718,
  154, 167, 156, 719,
  155, 168, 289, 720,
  24, 169, 158, 145,
  157, 170, 159, 146,
  158, 171, 160, 147,
  159, 172, 161, 148,
  160, 173, 162, 149,
  161, 174, 163, 150,
  162, 175, 164, 151,
  163, 176, 165, 152,
  164, 177, 166, 153,
  165, 178, 167, 154,
  166, 179, 168, 155,
  167, 180, 301, 156,
  36, 181, 170, 157,
  169, 182, 171, 158,
  170, 183, 172, 159,
  171, 184, 173, 160,
  172, 185, 174, 161,
  173, 186, 175, 162,
  174, 187, 176, 163,
  175, 188, 177, 164,
  176, 189, 178, 165,
  177, 190, 179, 166,
  178, 191, 180, 167,
  179, 192, 313, 168,
  48, 193, 182, 169,
  181, 194, 183, 170,
  182, 195, 184, 171,
  183, 196, 185, 172,
  184, 197, 186, 173,
  185, 198, 187, 174,
  186, 199, 188, 175,
  187, 200, 189, 176,
  188, 201, 190, 177,
  189, 202, 191, 178,
  190, 203, 192, 179,
  191, 204, 325, 180,
  60, 205, 194, 181,
  193, 206, 195, 182,
  194, 207, 196, 183,
  195, 208, 197, 184,
  196, 209, 198, 185,
  197, 210, 199, 186,
  198, 211, 200, 187,
  199, 212, 201, 188,
  200, 213, 202, 189,
  201, 214, 203, 190,
  202, 215, 204, 191,
  203, 216, 337, 192,
  72, 217, 206, 193,
  205, 218, 207, 194,
  206, 219, 208, 195,
  207, 220, 209, 196,
  208, 221, 210, 197,
  209, 222, 211, 198,
  210, 223, 212, 199,
  211, 224, 213, 200,
  212, 225, 214, 201,
  213, 226, 215, 202,
  214, 227, 216, 203,
  215, 228, 349, 204,
  84, 229, 218, 205,
  217, 230, 219, 206,
  218, 231, 220, 207,
  219, 232, 221, 208,
  220, 233, 222, 209,
  221, 234, 223, 210,
  222, 235, 224, 211,
  223, 236, 225, 212,
  224, 237, 226, 213,
  225, 238, 227, 214,
  226, 239, 228, 215,
  227, 240, 361, 216,
  96, 241, 230, 217,
  229, 242, 231, 218,
  230, 243, 232, 219,
  231, 244, 233, 220,
  232, 245, 234, 221,
  233, 246, 235, 222,
  234, 247, 236, 223,
  235, 248, 237, 224,
  236, 249, 238, 225,
  237, 250, 239, 226,
  238, 251, 240, 227,
  239, 252, 373, 228,
  108, 253, 242, 229,
  241, 254, 243, 230,
  242, 255, 244, 231,
  243, 256, 245, 232,
  244, 257, 246, 233,
  245, 258, 247, 234,
  246, 259, 248, 235,
  247, 260, 249, 236,
  248, 261, 250, 237,
  249, 262, 251, 238,
  250, 263, 252, 239,
  251, 264, 385, 240,
  120, 265, 254, 241,
  253, 266, 255, 242,
  254, 267, 256, 243,
  255, 268, 257, 244,
  256, 269, 258, 245,
  257, 270, 259, 246,
  258, 271, 260, 247,
  259, 272, 261, 248,
  260, 273, 262, 249,
  261, 274, 263, 250,
  262, 275, 264, 251,
  263, 276, 397, 252,
  132, 277, 266, 253,
  265, 278, 267, 254,
  266, 279, 268, 255,
  267, 280, 269, 256,
  268, 281, 270, 257,
  269, 282, 271, 258,
  270, 283, 272, 259,
  271, 284, 273, 260,
  272, 285, 274, 261,
  273, 286, 275, 262,
  274, 287, 276, 263,
  275, 288, 409, 264,
  144, 721, 278, 265,
  277, 722, 279, 266,
  278, 723, 280, 267,
  279, 724, 281, 268,
  280, 725, 282, 269,
  281, 726, 283, 270,
  282, 727, 284, 271,
  283, 728, 285, 272,
  284, 729, 286, 273,
  285, 730, 287, 274,
  286, 731, 288, 275,
  287, 732, 421, 276,
  301, 290, 720, 156,
  302, 291, 708, 289,
  303, 292, 696, 290,
  304, 293, 684, 291,
  305, 294, 672, 292,
  306, 295, 660, 293,
  307, 296, 648, 294,
  308, 297, 636, 295,
  309, 298, 624, 296,
  310, 299, 612, 297,
  311, 300, 600, 298,
  312, 433, 588, 299,
  313, 302, 289, 168,
  314, 303, 290, 301,
  315, 304, 291, 302,
  316, 305, 292, 303,
  317, 306, 293, 304,
  318, 307, 294, 305,
  319, 308, 295, 306,
  320, 309, 296, 307,
  321, 310, 297, 308,
  322, 311, 298, 309,
  323, 312, 299, 310,
  324, 445, 300, 311,
  325, 314, 301, 180,
  326, 315, 302, 313,
  327, 316, 303, 314,
  328, 317, 304, 315,
  329, 318, 305, 316,
  330, 319, 306, 317,
  331, 320, 307, 318,
  332, 321, 308, 319,
  333, 322, 309, 320,
  334, 323, 310, 321,
  335, 324, 311, 322,
  336, 457, 312, 323,
  337, 326, 313, 192,
  338, 327, 314, 325,
  339, 328, 315, 326,
  340, 329, 316, 327,
  341, 330, 317, 328,
  342, 331, 318, 329,
  343, 332, 319, 330,
  344, 333, 320, 331,
  345, 334, 321, 332,
  346, 335, 322, 333,
  347, 336, 323, 334,
  348, 469, 324, 335,
  349, 338, 325, 204,
  350, 339, 326, 337,
  351, 340, 327, 338,
  352, 341, 328, 339,
  353, 342, 329, 340,
  354, 343, 330, 341,
  355, 344, 331, 342,
  356, 345, 332, 343,
  357, 346, 333, 344,
  358, 347, 334, 345,
  359, 348, 335, 346,
  360, 481, 336, 347,
  361, 350, 337, 216,
  362, 351, 338, 349,
  363, 352, 339, 350,
  364, 353, 340, 351,
  365, 354, 341, 352,
  366, 355, 342, 353,
  367, 356, 343, 354,
  368, 357, 344, 355,
  369, 358, 345, 356,
  370, 359, 346, 357,
  371, 360, 347, 358,
  372, 493, 348, 359,
  373, 362, 349, 228,
  374, 363, 350, 361,
  375, 364, 351, 362,
  376, 365, 352, 363,
  377, 366, 353, 364,
  378, 367, 354, 365,
  379, 368, 355, 366,
  380, 369, 356, 367,
  381, 370, 357, 368,
  382, 371, 358, 369,
  383, 372, 359, 370,
  384, 505, 360, 371,
  385, 374, 361, 240,
  386, 375, 362, 373,
  387, 376, 363, 374,
  388, 377, 364, 375,
  389, 378, 365, 376,
  390, 379, 366, 377,
  391, 380, 367, 378,
  392, 381, 368, 379,
  393, 382, 369, 380,
  394, 383, 370, 381,
  395, 384, 371, 382,
  396, 517, 372, 383,
  397, 386, 373, 252,
  398, 387, 374, 385,
  399, 388, 375, 386,
  400, 389, 376, 387,
  401, 390, 377, 388,
  402, 391, 378, 389,
  403, 392, 379, 390,
  404, 393, 380, 391,
  405, 394, 381, 392,
  406, 395, 382, 393,
  407, 396, 383, 394,
  408, 529, 384, 395,
  409, 398, 385, 264,
  410, 399, 386, 397,
  411, 400, 387, 398,
  412, 401, 388, 399,
  413, 402, 389, 400,
  414, 403, 390, 401,
  415, 404, 391, 402,
  416, 405, 392, 403,
  417, 406, 393, 404,
  418, 407, 394, 405,
  419, 408, 395, 406,
  420, 541, 396, 407,
  421, 410, 397, 276,
  422, 411, 398, 409,
  423, 412, 399, 410,
  424, 413, 400, 411,
  425, 414, 401, 412,
  426, 415, 402, 413,
  427, 416, 403, 414,
  428, 417, 404, 415,
  429, 418, 405, 416,
  430, 419, 406, 417,
  431, 420, 407, 418,
  432, 553, 408, 419,
  732, 422, 409, 288,
  744, 423, 410, 421,
  756, 424, 411, 422,
  768, 425, 412, 423,
  780, 426, 413, 424,
  792, 427, 414, 425,
  804, 428, 415, 426,
  816, 429, 416, 427,
  828, 430, 417, 428,
  840, 431, 418, 429,
  852, 432, 419, 430,
  864, 565, 420, 431,
  445, 434, 588, 300,
  446, 435, 587, 433,
  447, 436, 586, 434,
  448, 437, 585, 435,
  449, 438, 584, 436,
  450, 439, 583, 437,
  451, 440, 582, 438,
  452, 441, 581, 439,
  453, 442, 580, 440,
  454, 443, 579, 441,
  455, 444, 578, 442,
  456, 1, 577, 443,
  457, 446, 433, 312,
  458, 447, 434, 445,
  459, 448, 435, 446,
  460, 449, 436, 447,
  461, 450, 437, 448,
  462, 451, 438, 449,
  463, 452, 439, 450,
  464, 453, 440, 451,
  465, 454, 441, 452,
  466, 455, 442, 453,
  467, 456, 443, 454,
  468, 13, 444, 455,
  469, 458, 445, 324,
  470, 459, 446, 457,
  471, 460, 447, 458,
  472, 461, 448, 459,
  473, 462, 449, 460,
  474, 463, 450, 461,
  475, 464, 451, 462,
  476, 465, 452, 463,
  477, 466, 453, 464,
  478, 467, 454, 465,
  479, 468, 455, 466,
  480, 25, 456, 467,
  481, 470, 457, 336,
  482, 471, 458, 469,
  483, 472, 459, 470,
  484, 473, 460, 471,
  485, 474, 461, 472,
  486, 475, 462, 473,
  487, 476, 463, 474,
  488, 477, 464, 475,
  489, 478, 465, 476,
  490, 479, 466, 477,
  491, 480, 467, 478,
  492, 37, 468, 479,
  493, 482, 469, 348,
  494, 483, 470, 481,
  495, 484, 471, 482,
  496, 485, 472, 483,
  497, 486, 473, 484,
  498, 487, 474, 485,
  499, 488, 475, 486,
  500, 489, 476, 487,
  501, 490, 477, 488,
  502, 491, 478, 489,
  503, 492, 479, 490,
  504, 49, 480, 491,
  505, 494, 481, 360,
  506, 495, 482, 493,
  507, 496, 483, 494,
  508, 497, 484, 495,
  509, 498, 485, 496,
  510, 499, 486, 497,
  511, 500, 487, 498,
  512, 501, 488, 499,
  513, 502, 489, 500,
  514, 503, 490, 501,
  515, 504, 491, 502,
  516, 61, 492, 503,
  517, 506, 493, 372,
  518, 507, 494, 505,
  519, 508, 495, 506,
  520, 509, 496, 507,
  521, 510, 497, 508,
  522, 511, 498, 509,
  523, 512, 499, 510,
  524, 513, 500, 511,
  525, 514, 501, 512,
  526, 515, 502, 513,
  527, 516, 503, 514,
  528, 73, 504, 515,
  529, 518, 505, 384,
  530, 519, 506, 517,
  531, 520, 507, 518,
  532, 521, 508, 519,
  533, 522, 509, 520,
  534, 523, 510, 521,
  535, 524, 511, 522,
  536, 525, 512, 523,
  537, 526, 513, 524,
  538, 527, 514, 525,
  539, 528, 515, 526,
  540, 85, 516, 527,
  541, 530, 517, 396,
  542, 531, 518, 529,
  543, 532, 519, 530,
  544, 533, 520, 531,
  545, 534, 521, 532,
  546, 535, 522, 533,
  547, 536, 523, 534,
  548, 537, 524, 535,
  549, 538, 525, 536,
  550, 539, 526, 537,
  551, 540, 527, 538,
  552, 97, 528, 539,
  553, 542, 529, 408,
  554, 543, 530, 541,
  555, 544, 531, 542,
  556, 545, 532, 543,
  557, 546, 533, 544,
  558, 547, 534, 545,
  559, 548, 535, 546,
  560, 549, 536, 547,
  561, 550, 537, 548,
  562, 551, 538, 549,
  563, 552, 539, 550,
  564, 109, 540, 551,
  565, 554, 541, 420,
  566, 555, 542, 553,
  567, 556, 543, 554,
  568, 557, 544, 555,
  569, 558, 545, 556,
  570, 559, 546, 557,
  571, 560, 547, 558,
  572, 561, 548, 559,
  573, 562, 549, 560,
  574, 563, 550, 561,
  575, 564, 551, 562,
  576, 121, 552, 563,
  864, 566, 553, 432,
  863, 567, 554, 565,
  862, 568, 555, 566,
  861, 569, 556, 567,
  860, 570, 557, 568,
  859, 571, 558, 569,
  858, 572, 559, 570,
  857, 573, 560, 571,
  856, 574, 561, 572,
  855, 575, 562, 573,
  854, 576, 563, 574,
  853, 133, 564, 575,
  444, 1, 589, 578,
  443, 577, 590, 579,
  442, 578, 591, 580,
  441, 579, 592, 581,
  440, 580, 593, 582,
  439, 581, 594, 583,
  438, 582, 595, 584,
  437, 583, 596, 585,
  436, 584, 597, 586,
  435, 585, 598, 587,
  434, 586, 599, 588,
  433, 587, 600, 300,
  577, 2, 601, 590,
  578, 589, 602, 591,
  579, 590, 603, 592,
  580, 591, 604, 593,
  581, 592, 605, 594,
  582, 593, 606, 595,
  583, 594, 607, 596,
  584, 595, 608, 597,
  585, 596, 609, 598,
  586, 597, 610, 599,
  587, 598, 611, 600,
  588, 599, 612, 299,
  589, 3, 613, 602,
  590, 601, 614, 603,
  591, 602, 615, 604,
  592, 603, 616, 605,
  593, 604, 617, 606,
  594, 605, 618, 607,
  595, 606, 619, 608,
  596, 607, 620, 609,
  597, 608, 621, 610,
  598, 609, 622, 611,
  599, 610, 623, 612,
  600, 611, 624, 298,
  601, 4, 625, 614,
  602, 613, 626, 615,
  603, 614, 627, 616,
  604, 615, 628, 617,
  605, 616, 629, 618,
  606, 617, 630, 619,
  607, 618, 631, 620,
  608, 619, 632, 621,
  609, 620, 633, 622,
  610, 621, 634, 623,
  611, 622, 635, 624,
  612, 623, 636, 297,
  613, 5, 637, 626,
  614, 625, 638, 627,
  615, 626, 639, 628,
  616, 627, 640, 629,
  617, 628, 641, 630,
  618, 629, 642, 631,
  619, 630, 643, 632,
  620, 631, 644, 633,
  621, 632, 645, 634,
  622, 633, 646, 635,
  623, 634, 647, 636,
  624, 635, 648, 296,
  625, 6, 649, 638,
  626, 637, 650, 639,
  627, 638, 651, 640,
  628, 639, 652, 641,
  629, 640, 653, 642,
  630, 641, 654, 643,
  631, 642, 655, 644,
  632, 643, 656, 645,
  633, 644, 657, 646,
  634, 645, 658, 647,
  635, 646, 659, 648,
  636, 647, 660, 295,
  637, 7, 661, 650,
  638, 649, 662, 651,
  639, 650, 663, 652,
  640, 651, 664, 653,
  641, 652, 665, 654,
  642, 653, 666, 655,
  643, 654, 667, 656,
  644, 655, 668, 657,
  645, 656, 669, 658,
  646, 657, 670, 659,
  647, 658, 671, 660,
  648, 659, 672, 294,
  649, 8, 673, 662,
  650, 661, 674, 663,
  651, 662, 675, 664,
  652, 663, 676, 665,
  653, 664, 677, 666,
  654, 665, 678, 667,
  655, 666, 679, 668,
  656, 667, 680, 669,
  657, 668, 681, 670,
  658, 669, 682, 671,
  659, 670, 683, 672,
  660, 671, 684, 293,
  661, 9, 685, 674,
  662, 673, 686, 675,
  663, 674, 687, 676,
  664, 675, 688, 677,
  665, 676, 689, 678,
  666, 677, 690, 679,
  667, 678, 691, 680,
  668, 679, 692, 681,
  669, 680, 693, 682,
  670, 681, 694, 683,
  671, 682, 695, 684,
  672, 683, 696, 292,
  673, 10, 697, 686,
  674, 685, 698, 687,
  675, 686, 699, 688,
  676, 687, 700, 689,
  677, 688, 701, 690,
  678, 689, 702, 691,
  679, 690, 703, 692,
  680, 691, 704, 693,
  681, 692, 705, 694,
  682, 693, 706, 695,
  683, 694, 707, 696,
  684, 695, 708, 291,
  685, 11, 709, 698,
  686, 697, 710, 699,
  687, 698, 711, 700,
  688, 699, 712, 701,
  689, 700, 713, 702,
  690, 701, 714, 703,
  691, 702, 715, 704,
  692, 703, 716, 705,
  693, 704, 717, 706,
  694, 705, 718, 707,
  695, 706, 719, 708,
  696, 707, 720, 290,
  697, 12, 145, 710,
  698, 709, 146, 711,
  699, 710, 147, 712,
  700, 711, 148, 713,
  701, 712, 149, 714,
  702, 713, 150, 715,
  703, 714, 151, 716,
  704, 715, 152, 717,
  705, 716, 153, 718,
  706, 717, 154, 719,
  707, 718, 155, 720,
  708, 719, 156, 289,
  144, 733, 722, 277,
  721, 734, 723, 278,
  722, 735, 724, 279,
  723, 736, 725, 280,
  724, 737, 726, 281,
  725, 738, 727, 282,
  726, 739, 728, 283,
  727, 740, 729, 284,
  728, 741, 730, 285,
  729, 742, 731, 286,
  730, 743, 732, 287,
  731, 744, 421, 288,
  143, 745, 734, 721,
  733, 746, 735, 722,
  734, 747, 736, 723,
  735, 748, 737, 724,
  736, 749, 738, 725,
  737, 750, 739, 726,
  738, 751, 740, 727,
  739, 752, 741, 728,
  740, 753, 742, 729,
  741, 754, 743, 730,
  742, 755, 744, 731,
  743, 756, 422, 732,
  142, 757, 746, 733,
  745, 758, 747, 734,
  746, 759, 748, 735,
  747, 760, 749, 736,
  748, 761, 750, 737,
  749, 762, 751, 738,
  750, 763, 752, 739,
  751, 764, 753, 740,
  752, 765, 754, 741,
  753, 766, 755, 742,
  754, 767, 756, 743,
  755, 768, 423, 744,
  141, 769, 758, 745,
  757, 770, 759, 746,
  758, 771, 760, 747,
  759, 772, 761, 748,
  760, 773, 762, 749,
  761, 774, 763, 750,
  762, 775, 764, 751,
  763, 776, 765, 752,
  764, 777, 766, 753,
  765, 778, 767, 754,
  766, 779, 768, 755,
  767, 780, 424, 756,
  140, 781, 770, 757,
  769, 782, 771, 758,
  770, 783, 772, 759,
  771, 784, 773, 760,
  772, 785, 774, 761,
  773, 786, 775, 762,
  774, 787, 776, 763,
  775, 788, 777, 764,
  776, 789, 778, 765,
  777, 790, 779, 766,
  778, 791, 780, 767,
  779, 792, 425, 768,
  139, 793, 782, 769,
  781, 794, 783, 770,
  782, 795, 784, 771,
  783, 796, 785, 772,
  784, 797, 786, 773,
  785, 798, 787, 774,
  786, 799, 788, 775,
  787, 800, 789, 776,
  788, 801, 790, 777,
  789, 802, 791, 778,
  790, 803, 792, 779,
  791, 804, 426, 780,
  138, 805, 794, 781,
  793, 806, 795, 782,
  794, 807, 796, 783,
  795, 808, 797, 784,
  796, 809, 798, 785,
  797, 810, 799, 786,
  798, 811, 800, 787,
  799, 812, 801, 788,
  800, 813, 802, 789,
  801, 814, 803, 790,
  802, 815, 804, 791,
  803, 816, 427, 792,
  137, 817, 806, 793,
  805, 818, 807, 794,
  806, 819, 808, 795,
  807, 820, 809, 796,
  808, 821, 810, 797,
  809, 822, 811, 798,
  810, 823, 812, 799,
  811, 824, 813, 800,
  812, 825, 814, 801,
  813, 826, 815, 802,
  814, 827, 816, 803,
  815, 828, 428, 804,
  136, 829, 818, 805,
  817, 830, 819, 806,
  818, 831, 820, 807,
  819, 832, 821, 808,
  820, 833, 822, 809,
  821, 834, 823, 810,
  822, 835, 824, 811,
  823, 836, 825, 812,
  824, 837, 826, 813,
  825, 838, 827, 814,
  826, 839, 828, 815,
  827, 840, 429, 816,
  135, 841, 830, 817,
  829, 842, 831, 818,
  830, 843, 832, 819,
  831, 844, 833, 820,
  832, 845, 834, 821,
  833, 846, 835, 822,
  834, 847, 836, 823,
  835, 848, 837, 824,
  836, 849, 838, 825,
  837, 850, 839, 826,
  838, 851, 840, 827,
  839, 852, 430, 828,
  134, 853, 842, 829,
  841, 854, 843, 830,
  842, 855, 844, 831,
  843, 856, 845, 832,
  844, 857, 846, 833,
  845, 858, 847, 834,
  846, 859, 848, 835,
  847, 860, 849, 836,
  848, 861, 850, 837,
  849, 862, 851, 838,
  850, 863, 852, 839,
  851, 864, 431, 840,
  133, 576, 854, 841,
  853, 575, 855, 842,
  854, 574, 856, 843,
  855, 573, 857, 844,
  856, 572, 858, 845,
  857, 571, 859, 846,
  858, 570, 860, 847,
  859, 569, 861, 848,
  860, 568, 862, 849,
  861, 567, 863, 850,
  862, 566, 864, 851,
  863, 565, 432, 852 ;

 dynamics_node_x = -45, -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 
    37.5, -45, -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, -45, 
    -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, -45, -37.5, 
    -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, -45, -37.5, -30, 
    -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, -45, -37.5, -30, -22.5, 
    -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, -45, -37.5, -30, -22.5, -15, -7.5, 
    0, 7.5, 15, 22.5, 30, 37.5, -45, -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 
    15, 22.5, 30, 37.5, -45, -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 
    30, 37.5, -45, -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, 
    -45, -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, -45, 
    -37.5, -30, -22.5, -15, -7.5, 0, 7.5, 15, 22.5, 30, 37.5, 45, 52.5, 60, 
    67.5, 75, 82.5, 90, 97.5, 105, 112.5, 120, 127.5, 45, 52.5, 60, 67.5, 75, 
    82.5, 90, 97.5, 105, 112.5, 120, 127.5, 45, 52.5, 60, 67.5, 75, 82.5, 90, 
    97.5, 105, 112.5, 120, 127.5, 45, 52.5, 60, 67.5, 75, 82.5, 90, 97.5, 
    105, 112.5, 120, 127.5, 45, 52.5, 60, 67.5, 75, 82.5, 90, 97.5, 105, 
    112.5, 120, 127.5, 45, 52.5, 60, 67.5, 75, 82.5, 90, 97.5, 105, 112.5, 
    120, 127.5, 45, 52.5, 60, 67.5, 75, 82.5, 90, 97.5, 105, 112.5, 120, 
    127.5, 45, 52.5, 60, 67.5, 75, 82.5, 90, 97.5, 105, 112.5, 120, 127.5, 
    45, 52.5, 60, 67.5, 75, 82.5, 90, 97.5, 105, 112.5, 120, 127.5, 45, 52.5, 
    60, 67.5, 75, 82.5, 90, 97.5, 105, 112.5, 120, 127.5, 45, 52.5, 60, 67.5, 
    75, 82.5, 90, 97.5, 105, 112.5, 120, 127.5, 45, 52.5, 60, 67.5, 75, 82.5, 
    90, 97.5, 105, 112.5, 120, 127.5, 135, 142.5, 150, 157.5, 165, 172.5, 
    -180, -172.5, -165, -157.5, -150, -142.5, 135, 142.5, 150, 157.5, 165, 
    172.5, -180, -172.5, -165, -157.5, -150, -142.5, 135, 142.5, 150, 157.5, 
    165, 172.5, -180, -172.5, -165, -157.5, -150, -142.5, 135, 142.5, 150, 
    157.5, 165, 172.5, -180, -172.5, -165, -157.5, -150, -142.5, 135, 142.5, 
    150, 157.5, 165, 172.5, -180, -172.5, -165, -157.5, -150, -142.5, 135, 
    142.5, 150, 157.5, 165, 172.5, -180, -172.5, -165, -157.5, -150, -142.5, 
    135, 142.5, 150, 157.5, 165, 172.5, -180, -172.5, -165, -157.5, -150, 
    -142.5, 135, 142.5, 150, 157.5, 165, 172.5, -180, -172.5, -165, -157.5, 
    -150, -142.5, 135, 142.5, 150, 157.5, 165, 172.5, -180, -172.5, -165, 
    -157.5, -150, -142.5, 135, 142.5, 150, 157.5, 165, 172.5, -180, -172.5, 
    -165, -157.5, -150, -142.5, 135, 142.5, 150, 157.5, 165, 172.5, -180, 
    -172.5, -165, -157.5, -150, -142.5, 135, 142.5, 150, 157.5, 165, 172.5, 
    -180, -172.5, -165, -157.5, -150, -142.5, -135, -127.5, -120, -112.5, 
    -105, -97.5, -90, -82.5, -75, -67.5, -60, -52.5, -135, -127.5, -120, 
    -112.5, -105, -97.5, -90, -82.5, -75, -67.5, -60, -52.5, -135, -127.5, 
    -120, -112.5, -105, -97.5, -90, -82.5, -75, -67.5, -60, -52.5, -135, 
    -127.5, -120, -112.5, -105, -97.5, -90, -82.5, -75, -67.5, -60, -52.5, 
    -135, -127.5, -120, -112.5, -105, -97.5, -90, -82.5, -75, -67.5, -60, 
    -52.5, -135, -127.5, -120, -112.5, -105, -97.5, -90, -82.5, -75, -67.5, 
    -60, -52.5, -135, -127.5, -120, -112.5, -105, -97.5, -90, -82.5, -75, 
    -67.5, -60, -52.5, -135, -127.5, -120, -112.5, -105, -97.5, -90, -82.5, 
    -75, -67.5, -60, -52.5, -135, -127.5, -120, -112.5, -105, -97.5, -90, 
    -82.5, -75, -67.5, -60, -52.5, -135, -127.5, -120, -112.5, -105, -97.5, 
    -90, -82.5, -75, -67.5, -60, -52.5, -135, -127.5, -120, -112.5, -105, 
    -97.5, -90, -82.5, -75, -67.5, -60, -52.5, -135, -127.5, -120, -112.5, 
    -105, -97.5, -90, -82.5, -75, -67.5, -60, -52.5, -45, -53.04155641726, 
    -61.6392220370136, -70.7508909984478, -80.2643896827547, -90, 
    -99.7356103172453, -109.249109001552, -118.360777962986, 
    -126.95844358274, -135, -36.95844358274, -45, -54.3428701752672, 
    -65.1039093610171, -77.1545477812505, -90, -102.84545221875, 
    -114.896090638983, -125.657129824733, -135, -143.04155641726, 
    -28.3607779629864, -35.6571298247328, -45, -57.1017141696649, 
    -72.3678051586227, -90, -107.632194841377, -122.898285830335, -135, 
    -144.342870175267, -151.639222037014, -19.2491090015522, 
    -24.8960906389829, -32.8982858303351, -45, -63.8335530583408, -90, 
    -116.166446941659, -135, -147.101714169665, -155.103909361017, 
    -160.750890998448, -9.73561031724535, -12.8454522187495, 
    -17.6321948413773, -26.1664469416592, -45, -90, -135, -153.833553058341, 
    -162.367805158623, -167.15454778125, -170.264389682755, 0, 0, 0, 0, 0, 0, 
    -180, -180, -180, -180, -180, 9.73561031724534, 12.8454522187495, 
    17.6321948413773, 26.1664469416592, 45, 90, 135, 153.833553058341, 
    162.367805158623, 167.15454778125, 170.264389682755, 19.2491090015522, 
    24.8960906389829, 32.8982858303351, 45, 63.8335530583408, 90, 
    116.166446941659, 135, 147.101714169665, 155.103909361017, 
    160.750890998448, 28.3607779629864, 35.6571298247328, 45, 
    57.1017141696649, 72.3678051586227, 90, 107.632194841377, 
    122.898285830335, 135, 144.342870175267, 151.639222037014, 
    36.95844358274, 45, 54.3428701752672, 65.1039093610171, 77.1545477812505, 
    90, 102.84545221875, 114.896090638983, 125.657129824733, 135, 
    143.04155641726, 45, 53.0415564172599, 61.6392220370136, 
    70.7508909984478, 80.2643896827547, 90, 99.7356103172453, 
    109.249109001552, 118.360777962986, 126.95844358274, 135, 45, 52.5, 60, 
    67.5, 75, 82.5, 90, 97.5, 105, 112.5, 120, 127.5, 37.5, 45, 
    53.04155641726, 61.6392220370136, 70.7508909984478, 80.2643896827547, 90, 
    99.7356103172453, 109.249109001552, 118.360777962986, 126.95844358274, 
    135, 30, 36.95844358274, 45, 54.3428701752672, 65.1039093610171, 
    77.1545477812505, 90, 102.84545221875, 114.896090638983, 
    125.657129824733, 135, 143.04155641726, 22.5, 28.3607779629864, 
    35.6571298247328, 45, 57.1017141696649, 72.3678051586227, 90, 
    107.632194841377, 122.898285830335, 135, 144.342870175267, 
    151.639222037014, 15, 19.2491090015522, 24.8960906389829, 
    32.8982858303351, 45, 63.8335530583408, 90, 116.166446941659, 135, 
    147.101714169665, 155.103909361017, 160.750890998448, 7.50000000000001, 
    9.73561031724535, 12.8454522187495, 17.6321948413773, 26.1664469416592, 
    45, 90, 135, 153.833553058341, 162.367805158623, 167.15454778125, 
    170.264389682755, -0, -0, -0, -0, -0, -0, 0, -180, -180, -180, -180, 
    -180, -7.5, -9.73561031724534, -12.8454522187495, -17.6321948413773, 
    -26.1664469416592, -45, -90, -135, -153.833553058341, -162.367805158623, 
    -167.15454778125, -170.264389682755, -15, -19.2491090015522, 
    -24.8960906389829, -32.8982858303351, -45, -63.8335530583408, -90, 
    -116.166446941659, -135, -147.101714169665, -155.103909361017, 
    -160.750890998448, -22.5, -28.3607779629864, -35.6571298247328, -45, 
    -57.1017141696649, -72.3678051586227, -90, -107.632194841377, 
    -122.898285830335, -135, -144.342870175267, -151.639222037014, -30, 
    -36.95844358274, -45, -54.3428701752672, -65.1039093610171, 
    -77.1545477812505, -90, -102.84545221875, -114.896090638983, 
    -125.657129824733, -135, -143.04155641726, -37.5, -45, -53.0415564172599, 
    -61.6392220370136, -70.7508909984478, -80.2643896827547, -90, 
    -99.7356103172453, -109.249109001552, -118.360777962986, 
    -126.95844358274, -135, -45, -52.5, -60, -67.5, -75, -82.5, -90, -97.5, 
    -105, -112.5, -120, -127.5, 135, 142.5, 150, 157.5, 165, 172.5, -180, 
    -172.5, -165, -157.5, -150, -142.5, -135 ;

 dynamics_node_y = 35.2643896827547, 38.4268434976953, 40.8933946491309, 
    42.7342096008998, 44.0070271956363, 44.753861966975, 45, 44.753861966975, 
    44.0070271956363, 42.7342096008998, 40.8933946491309, 38.4268434976953, 
    28.4834661179317, 31.3314426644734, 33.6050181915629, 35.3335026120138, 
    36.5451381553822, 37.2625128714784, 37.5, 37.2625128714784, 
    36.5451381553822, 35.3335026120138, 33.6050181915629, 31.3314426644734, 
    22.2076542985965, 24.6098050837908, 26.565051177078, 28.0755542102809, 
    29.1474262640282, 29.7872947635816, 30, 29.7872947635816, 
    29.1474262640282, 28.0755542102809, 26.565051177078, 24.6098050837908, 
    16.3249499368952, 18.1914391843494, 19.7338984646069, 20.9410204722438, 
    21.8063277400641, 22.3264806874313, 22.5, 22.3264806874313, 
    21.8063277400641, 20.9410204722438, 19.7338984646069, 18.1914391843494, 
    10.7285831216091, 12.0011964297362, 13.0643134295083, 13.9041999653766, 
    14.5108186990699, 14.8773865849752, 15, 14.8773865849752, 
    14.5108186990699, 13.9041999653766, 13.0643134295083, 12.0011964297362, 
    5.31847183939939, 5.96274919276321, 6.50445695752584, 6.93488111564006, 
    7.247207855436, 7.43655768147728, 7.5, 7.43655768147728, 7.247207855436, 
    6.93488111564006, 6.50445695752584, 5.96274919276321, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -5.31847183939939, -5.9627491927632, 
    -6.50445695752584, -6.93488111564005, -7.24720785543599, 
    -7.43655768147727, -7.5, -7.43655768147727, -7.24720785543599, 
    -6.93488111564005, -6.50445695752584, -5.9627491927632, 
    -10.7285831216091, -12.0011964297362, -13.0643134295083, 
    -13.9041999653766, -14.5108186990699, -14.8773865849752, -15, 
    -14.8773865849752, -14.5108186990699, -13.9041999653766, 
    -13.0643134295083, -12.0011964297362, -16.3249499368952, 
    -18.1914391843494, -19.7338984646069, -20.9410204722438, 
    -21.8063277400641, -22.3264806874313, -22.5, -22.3264806874313, 
    -21.8063277400641, -20.9410204722438, -19.7338984646069, 
    -18.1914391843494, -22.2076542985965, -24.6098050837908, 
    -26.565051177078, -28.0755542102809, -29.1474262640282, 
    -29.7872947635816, -30, -29.7872947635816, -29.1474262640282, 
    -28.0755542102809, -26.565051177078, -24.6098050837908, 
    -28.4834661179317, -31.3314426644734, -33.6050181915629, 
    -35.3335026120138, -36.5451381553822, -37.2625128714784, -37.5, 
    -37.2625128714784, -36.5451381553822, -35.3335026120138, 
    -33.6050181915629, -31.3314426644734, 35.2643896827547, 38.4268434976953, 
    40.8933946491309, 42.7342096008998, 44.0070271956363, 44.753861966975, 
    45, 44.753861966975, 44.0070271956363, 42.7342096008998, 
    40.8933946491309, 38.4268434976953, 28.4834661179317, 31.3314426644734, 
    33.6050181915629, 35.3335026120138, 36.5451381553822, 37.2625128714784, 
    37.5, 37.2625128714784, 36.5451381553822, 35.3335026120138, 
    33.6050181915629, 31.3314426644734, 22.2076542985965, 24.6098050837908, 
    26.565051177078, 28.0755542102809, 29.1474262640282, 29.7872947635816, 
    30, 29.7872947635816, 29.1474262640282, 28.0755542102809, 
    26.565051177078, 24.6098050837908, 16.3249499368952, 18.1914391843494, 
    19.7338984646069, 20.9410204722438, 21.8063277400641, 22.3264806874313, 
    22.5, 22.3264806874313, 21.8063277400641, 20.9410204722438, 
    19.7338984646069, 18.1914391843494, 10.7285831216091, 12.0011964297362, 
    13.0643134295083, 13.9041999653766, 14.5108186990699, 14.8773865849752, 
    15, 14.8773865849752, 14.5108186990699, 13.9041999653766, 
    13.0643134295083, 12.0011964297362, 5.31847183939939, 5.96274919276321, 
    6.50445695752584, 6.93488111564006, 7.247207855436, 7.43655768147728, 
    7.5, 7.43655768147728, 7.247207855436, 6.93488111564006, 
    6.50445695752584, 5.96274919276321, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -5.31847183939939, -5.9627491927632, -6.50445695752584, 
    -6.93488111564005, -7.24720785543599, -7.43655768147727, -7.5, 
    -7.43655768147727, -7.24720785543599, -6.93488111564005, 
    -6.50445695752584, -5.9627491927632, -10.7285831216091, 
    -12.0011964297362, -13.0643134295083, -13.9041999653766, 
    -14.5108186990699, -14.8773865849752, -15, -14.8773865849752, 
    -14.5108186990699, -13.9041999653766, -13.0643134295083, 
    -12.0011964297362, -16.3249499368952, -18.1914391843494, 
    -19.7338984646069, -20.9410204722438, -21.8063277400641, 
    -22.3264806874313, -22.5, -22.3264806874313, -21.8063277400641, 
    -20.9410204722438, -19.7338984646069, -18.1914391843494, 
    -22.2076542985965, -24.6098050837908, -26.565051177078, 
    -28.0755542102809, -29.1474262640282, -29.7872947635816, -30, 
    -29.7872947635816, -29.1474262640282, -28.0755542102809, 
    -26.565051177078, -24.6098050837908, -28.4834661179317, 
    -31.3314426644734, -33.6050181915629, -35.3335026120138, 
    -36.5451381553822, -37.2625128714784, -37.5, -37.2625128714784, 
    -36.5451381553822, -35.3335026120138, -33.6050181915629, 
    -31.3314426644734, 35.2643896827547, 38.4268434976953, 40.8933946491309, 
    42.7342096008998, 44.0070271956363, 44.753861966975, 45, 44.753861966975, 
    44.0070271956363, 42.7342096008998, 40.8933946491309, 38.4268434976953, 
    28.4834661179317, 31.3314426644734, 33.6050181915629, 35.3335026120138, 
    36.5451381553822, 37.2625128714784, 37.5, 37.2625128714784, 
    36.5451381553822, 35.3335026120138, 33.6050181915629, 31.3314426644734, 
    22.2076542985965, 24.6098050837908, 26.565051177078, 28.0755542102809, 
    29.1474262640282, 29.7872947635816, 30, 29.7872947635816, 
    29.1474262640282, 28.0755542102809, 26.565051177078, 24.6098050837908, 
    16.3249499368952, 18.1914391843494, 19.7338984646069, 20.9410204722438, 
    21.8063277400641, 22.3264806874313, 22.5, 22.3264806874313, 
    21.8063277400641, 20.9410204722438, 19.7338984646069, 18.1914391843494, 
    10.7285831216091, 12.0011964297362, 13.0643134295083, 13.9041999653766, 
    14.5108186990699, 14.8773865849752, 15, 14.8773865849752, 
    14.5108186990699, 13.9041999653766, 13.0643134295083, 12.0011964297362, 
    5.31847183939939, 5.96274919276321, 6.50445695752584, 6.93488111564006, 
    7.247207855436, 7.43655768147728, 7.5, 7.43655768147728, 7.247207855436, 
    6.93488111564006, 6.50445695752584, 5.96274919276321, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -5.31847183939939, -5.9627491927632, 
    -6.50445695752584, -6.93488111564005, -7.24720785543599, 
    -7.43655768147727, -7.5, -7.43655768147727, -7.24720785543599, 
    -6.93488111564005, -6.50445695752584, -5.9627491927632, 
    -10.7285831216091, -12.0011964297362, -13.0643134295083, 
    -13.9041999653766, -14.5108186990699, -14.8773865849752, -15, 
    -14.8773865849752, -14.5108186990699, -13.9041999653766, 
    -13.0643134295083, -12.0011964297362, -16.3249499368952, 
    -18.1914391843494, -19.7338984646069, -20.9410204722438, 
    -21.8063277400641, -22.3264806874313, -22.5, -22.3264806874313, 
    -21.8063277400641, -20.9410204722438, -19.7338984646069, 
    -18.1914391843494, -22.2076542985965, -24.6098050837908, 
    -26.565051177078, -28.0755542102809, -29.1474262640282, 
    -29.7872947635816, -30, -29.7872947635816, -29.1474262640282, 
    -28.0755542102809, -26.565051177078, -24.6098050837908, 
    -28.4834661179317, -31.3314426644734, -33.6050181915629, 
    -35.3335026120138, -36.5451381553822, -37.2625128714784, -37.5, 
    -37.2625128714784, -36.5451381553822, -35.3335026120138, 
    -33.6050181915629, -31.3314426644734, 35.2643896827547, 38.4268434976953, 
    40.8933946491309, 42.7342096008998, 44.0070271956363, 44.753861966975, 
    45, 44.753861966975, 44.0070271956363, 42.7342096008998, 
    40.8933946491309, 38.4268434976953, 28.4834661179317, 31.3314426644734, 
    33.6050181915629, 35.3335026120138, 36.5451381553822, 37.2625128714784, 
    37.5, 37.2625128714784, 36.5451381553822, 35.3335026120138, 
    33.6050181915629, 31.3314426644734, 22.2076542985965, 24.6098050837908, 
    26.565051177078, 28.0755542102809, 29.1474262640282, 29.7872947635816, 
    30, 29.7872947635816, 29.1474262640282, 28.0755542102809, 
    26.565051177078, 24.6098050837908, 16.3249499368952, 18.1914391843494, 
    19.7338984646069, 20.9410204722438, 21.8063277400641, 22.3264806874313, 
    22.5, 22.3264806874313, 21.8063277400641, 20.9410204722438, 
    19.7338984646069, 18.1914391843494, 10.7285831216091, 12.0011964297362, 
    13.0643134295083, 13.9041999653766, 14.5108186990699, 14.8773865849752, 
    15, 14.8773865849752, 14.5108186990699, 13.9041999653766, 
    13.0643134295083, 12.0011964297362, 5.31847183939939, 5.96274919276321, 
    6.50445695752584, 6.93488111564006, 7.247207855436, 7.43655768147728, 
    7.5, 7.43655768147728, 7.247207855436, 6.93488111564006, 
    6.50445695752584, 5.96274919276321, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -5.31847183939939, -5.9627491927632, -6.50445695752584, 
    -6.93488111564005, -7.24720785543599, -7.43655768147727, -7.5, 
    -7.43655768147727, -7.24720785543599, -6.93488111564005, 
    -6.50445695752584, -5.9627491927632, -10.7285831216091, 
    -12.0011964297362, -13.0643134295083, -13.9041999653766, 
    -14.5108186990699, -14.8773865849752, -15, -14.8773865849752, 
    -14.5108186990699, -13.9041999653766, -13.0643134295083, 
    -12.0011964297362, -16.3249499368952, -18.1914391843494, 
    -19.7338984646069, -20.9410204722438, -21.8063277400641, 
    -22.3264806874313, -22.5, -22.3264806874313, -21.8063277400641, 
    -20.9410204722438, -19.7338984646069, -18.1914391843494, 
    -22.2076542985965, -24.6098050837908, -26.565051177078, 
    -28.0755542102809, -29.1474262640282, -29.7872947635816, -30, 
    -29.7872947635816, -29.1474262640282, -28.0755542102809, 
    -26.565051177078, -24.6098050837908, -28.4834661179317, 
    -31.3314426644734, -33.6050181915629, -35.3335026120138, 
    -36.5451381553822, -37.2625128714784, -37.5, -37.2625128714784, 
    -36.5451381553822, -35.3335026120138, -33.6050181915629, 
    -31.3314426644734, 42.6611719623651, 46.1610034997872, 48.9119528722244, 
    50.8969852747691, 52.0978484161962, 52.5, 52.0978484161962, 
    50.8969852747691, 48.9119528722244, 46.1610034997872, 42.6611719623651, 
    46.1610034997872, 50.7684795164077, 54.6036351534441, 57.5233157615547, 
    59.3672407834663, 60, 59.3672407834663, 57.5233157615547, 
    54.6036351534441, 50.7684795164078, 46.1610034997872, 48.9119528722244, 
    54.6036351534441, 59.6388065951783, 63.7417202794995, 66.5086765471698, 
    67.5, 66.5086765471698, 63.7417202794995, 59.6388065951783, 
    54.6036351534441, 48.9119528722244, 50.8969852747691, 57.5233157615547, 
    63.7417202794995, 69.2464290163152, 73.3772654499124, 75, 
    73.3772654499124, 69.2464290163152, 63.7417202794995, 57.5233157615548, 
    50.8969852747691, 52.0978484161962, 59.3672407834663, 66.5086765471698, 
    73.3772654499124, 79.453161100789, 82.5, 79.453161100789, 
    73.3772654499124, 66.5086765471698, 59.3672407834663, 52.0978484161962, 
    52.5, 60, 67.5, 75, 82.5, 90, 82.5, 75, 67.5, 60, 52.5, 52.0978484161962, 
    59.3672407834663, 66.5086765471698, 73.3772654499124, 79.453161100789, 
    82.5, 79.453161100789, 73.3772654499124, 66.5086765471698, 
    59.3672407834663, 52.0978484161962, 50.8969852747691, 57.5233157615547, 
    63.7417202794995, 69.2464290163152, 73.3772654499124, 75, 
    73.3772654499124, 69.2464290163152, 63.7417202794995, 57.5233157615548, 
    50.8969852747691, 48.9119528722244, 54.6036351534441, 59.6388065951783, 
    63.7417202794995, 66.5086765471698, 67.5, 66.5086765471698, 
    63.7417202794995, 59.6388065951783, 54.6036351534441, 48.9119528722244, 
    46.1610034997872, 50.7684795164078, 54.6036351534441, 57.5233157615548, 
    59.3672407834663, 60, 59.3672407834663, 57.5233157615548, 
    54.6036351534441, 50.7684795164078, 46.1610034997873, 42.6611719623651, 
    46.1610034997872, 48.9119528722244, 50.8969852747691, 52.0978484161962, 
    52.5, 52.0978484161962, 50.8969852747691, 48.9119528722244, 
    46.1610034997873, 42.6611719623651, -35.2643896827547, -38.4268434976953, 
    -40.8933946491309, -42.7342096008998, -44.0070271956363, 
    -44.753861966975, -45, -44.753861966975, -44.0070271956363, 
    -42.7342096008998, -40.8933946491309, -38.4268434976953, 
    -38.4268434976953, -42.6611719623651, -46.1610034997872, 
    -48.9119528722244, -50.8969852747691, -52.0978484161962, -52.5, 
    -52.0978484161962, -50.8969852747691, -48.9119528722244, 
    -46.1610034997872, -42.6611719623651, -40.8933946491309, 
    -46.1610034997872, -50.7684795164077, -54.6036351534441, 
    -57.5233157615547, -59.3672407834663, -60, -59.3672407834663, 
    -57.5233157615547, -54.6036351534441, -50.7684795164078, 
    -46.1610034997872, -42.7342096008998, -48.9119528722244, 
    -54.6036351534441, -59.6388065951783, -63.7417202794995, 
    -66.5086765471698, -67.5, -66.5086765471698, -63.7417202794995, 
    -59.6388065951783, -54.6036351534441, -48.9119528722244, 
    -44.0070271956363, -50.8969852747691, -57.5233157615547, 
    -63.7417202794995, -69.2464290163152, -73.3772654499124, -75, 
    -73.3772654499124, -69.2464290163152, -63.7417202794995, 
    -57.5233157615548, -50.8969852747691, -44.753861966975, 
    -52.0978484161962, -59.3672407834663, -66.5086765471698, 
    -73.3772654499124, -79.453161100789, -82.5, -79.453161100789, 
    -73.3772654499124, -66.5086765471698, -59.3672407834663, 
    -52.0978484161962, -45, -52.5, -60, -67.5, -75, -82.5, -90, -82.5, -75, 
    -67.5, -60, -52.5, -44.753861966975, -52.0978484161962, 
    -59.3672407834663, -66.5086765471698, -73.3772654499124, 
    -79.453161100789, -82.5, -79.453161100789, -73.3772654499124, 
    -66.5086765471698, -59.3672407834663, -52.0978484161962, 
    -44.0070271956363, -50.8969852747691, -57.5233157615547, 
    -63.7417202794995, -69.2464290163152, -73.3772654499124, -75, 
    -73.3772654499124, -69.2464290163152, -63.7417202794995, 
    -57.5233157615548, -50.8969852747691, -42.7342096008998, 
    -48.9119528722244, -54.6036351534441, -59.6388065951783, 
    -63.7417202794995, -66.5086765471698, -67.5, -66.5086765471698, 
    -63.7417202794995, -59.6388065951783, -54.6036351534441, 
    -48.9119528722244, -40.8933946491309, -46.1610034997872, 
    -50.7684795164078, -54.6036351534441, -57.5233157615548, 
    -59.3672407834663, -60, -59.3672407834663, -57.5233157615548, 
    -54.6036351534441, -50.7684795164078, -46.1610034997873, 
    -38.4268434976953, -42.6611719623651, -46.1610034997872, 
    -48.9119528722244, -50.8969852747691, -52.0978484161962, -52.5, 
    -52.0978484161962, -50.8969852747691, -48.9119528722244, 
    -46.1610034997873, -42.6611719623651, -35.2643896827547, 
    -38.4268434976953, -40.8933946491309, -42.7342096008998, 
    -44.0070271956363, -44.753861966975, -45, -44.753861966975, 
    -44.0070271956363, -42.7342096008998, -40.8933946491309, 
    -38.4268434976953, -35.2643896827547, -38.4268434976953, 
    -40.8933946491309, -42.7342096008998, -44.0070271956363, 
    -44.753861966975, -45, -44.753861966975, -44.0070271956363, 
    -42.7342096008998, -40.8933946491309, -38.4268434976953, -35.2643896827547 ;

 dynamics_face_x = -41.3152089030983, -33.806771088304, -26.2960492462929, 
    -18.7838104277648, -11.2706263664288, -3.75692946913451, 3.7569294691345, 
    11.2706263664288, 18.7838104277648, 26.2960492462929, 33.806771088304, 
    41.3152089030983, -41.2936109384805, -33.7887716035354, 
    -26.2819825548092, -18.7737791519095, -11.2646279062497, 
    -3.75493465965447, 3.75493465965447, 11.2646279062497, 18.7737791519095, 
    26.2819825548092, 33.7887716035354, 41.2936109384805, -41.2763945590034, 
    -33.773869868729, -26.2699713858559, -18.7650111229678, -11.259302201907, 
    -3.75314966175661, 3.75314966175661, 11.259302201907, 18.7650111229678, 
    26.2699713858559, 33.773869868729, 41.2763945590034, -41.2636238596043, 
    -33.7624809909733, -26.2605583606434, -18.7580048589284, 
    -11.2549899787732, -3.75169466260126, 3.75169466260126, 11.2549899787732, 
    18.7580048589284, 26.2605583606434, 33.7624809909732, 41.2636238596043, 
    -41.2552106377437, -33.7548156148214, -26.254105045772, 
    -18.7531312562048, -11.2519601891623, -3.7506671461934, 3.75066714619339, 
    11.2519601891623, 18.7531312562048, 26.254105045772, 33.7548156148213, 
    41.2552106377437, -41.2510401544502, -33.7509666749151, 
    -26.2508281137282, -18.7506341927028, -11.2503981200382, 
    -3.75013569437423, 3.75013569437423, 11.2503981200382, 18.7506341927028, 
    26.2508281137282, 33.7509666749151, 41.2510401544502, -41.2510401544502, 
    -33.7509666749151, -26.2508281137282, -18.7506341927028, 
    -11.2503981200382, -3.75013569437423, 3.75013569437423, 11.2503981200382, 
    18.7506341927028, 26.2508281137282, 33.7509666749151, 41.2510401544502, 
    -41.2552106377437, -33.7548156148214, -26.254105045772, 
    -18.7531312562048, -11.2519601891623, -3.7506671461934, 3.75066714619339, 
    11.2519601891623, 18.7531312562048, 26.254105045772, 33.7548156148213, 
    41.2552106377437, -41.2636238596043, -33.7624809909732, 
    -26.2605583606434, -18.7580048589284, -11.2549899787732, 
    -3.75169466260126, 3.75169466260126, 11.2549899787732, 18.7580048589284, 
    26.2605583606434, 33.7624809909732, 41.2636238596043, -41.2763945590034, 
    -33.773869868729, -26.2699713858559, -18.7650111229678, -11.259302201907, 
    -3.75314966175661, 3.75314966175661, 11.259302201907, 18.7650111229678, 
    26.2699713858559, 33.773869868729, 41.2763945590034, -41.2936109384805, 
    -33.7887716035354, -26.2819825548092, -18.7737791519095, 
    -11.2646279062497, -3.75493465965447, 3.75493465965447, 11.2646279062497, 
    18.7737791519095, 26.2819825548092, 33.7887716035353, 41.2936109384805, 
    -41.3152089030983, -33.806771088304, -26.2960492462929, 
    -18.7838104277648, -11.2706263664288, -3.75692946913451, 
    3.75692946913451, 11.2706263664288, 18.7838104277648, 26.2960492462929, 
    33.806771088304, 41.3152089030983, 48.6847910969017, 56.1932289116959, 
    63.7039507537071, 71.2161895722352, 78.7293736335712, 86.2430705308655, 
    93.7569294691345, 101.270626366429, 108.783810427765, 116.296049246293, 
    123.806771088304, 131.315208903098, 48.7063890615195, 56.2112283964646, 
    63.7180174451908, 71.2262208480905, 78.7353720937503, 86.2450653403455, 
    93.7549346596545, 101.26462790625, 108.773779151909, 116.281982554809, 
    123.788771603535, 131.293610938481, 48.7236054409966, 56.226130131271, 
    63.7300286141441, 71.2349888770322, 78.740697798093, 86.2468503382434, 
    93.7531496617566, 101.259302201907, 108.765011122968, 116.269971385856, 
    123.773869868729, 131.276394559003, 48.7363761403957, 56.2375190090268, 
    63.7394416393566, 71.2419951410716, 78.7450100212268, 86.2483053373987, 
    93.7516946626012, 101.254989978773, 108.758004858928, 116.260558360643, 
    123.762480990973, 131.263623859604, 48.7447893622563, 56.2451843851786, 
    63.745894954228, 71.2468687437952, 78.7480398108377, 86.2493328538066, 
    93.7506671461934, 101.251960189162, 108.753131256205, 116.254105045772, 
    123.754815614821, 131.255210637744, 48.7489598455498, 56.2490333250849, 
    63.7491718862718, 71.2493658072972, 78.7496018799618, 86.2498643056258, 
    93.7501356943742, 101.250398120038, 108.750634192703, 116.250828113728, 
    123.750966674915, 131.25104015445, 48.7489598455498, 56.2490333250849, 
    63.7491718862718, 71.2493658072972, 78.7496018799618, 86.2498643056258, 
    93.7501356943742, 101.250398120038, 108.750634192703, 116.250828113728, 
    123.750966674915, 131.25104015445, 48.7447893622563, 56.2451843851786, 
    63.745894954228, 71.2468687437952, 78.7480398108377, 86.2493328538066, 
    93.7506671461934, 101.251960189162, 108.753131256205, 116.254105045772, 
    123.754815614821, 131.255210637744, 48.7363761403957, 56.2375190090268, 
    63.7394416393566, 71.2419951410716, 78.7450100212268, 86.2483053373987, 
    93.7516946626012, 101.254989978773, 108.758004858928, 116.260558360643, 
    123.762480990973, 131.263623859604, 48.7236054409966, 56.226130131271, 
    63.7300286141441, 71.2349888770322, 78.740697798093, 86.2468503382434, 
    93.7531496617566, 101.259302201907, 108.765011122968, 116.269971385856, 
    123.773869868729, 131.276394559003, 48.7063890615195, 56.2112283964646, 
    63.7180174451908, 71.2262208480905, 78.7353720937503, 86.2450653403455, 
    93.7549346596545, 101.26462790625, 108.773779151909, 116.281982554809, 
    123.788771603535, 131.293610938481, 48.6847910969017, 56.193228911696, 
    63.7039507537071, 71.2161895722352, 78.7293736335712, 86.2430705308655, 
    93.7569294691345, 101.270626366429, 108.783810427765, 116.296049246293, 
    123.806771088304, 131.315208903098, 138.684791096902, 146.193228911696, 
    153.703950753707, 161.216189572235, 168.729373633571, 176.243070530866, 
    -176.243070530866, -168.729373633571, -161.216189572235, 
    -153.703950753707, -146.193228911696, -138.684791096902, 
    138.706389061519, 146.211228396465, 153.718017445191, 161.226220848091, 
    168.73537209375, 176.245065340346, -176.245065340346, -168.73537209375, 
    -161.226220848091, -153.718017445191, -146.211228396465, 
    -138.706389061519, 138.723605440997, 146.226130131271, 153.730028614144, 
    161.234988877032, 168.740697798093, 176.246850338243, -176.246850338243, 
    -168.740697798093, -161.234988877032, -153.730028614144, 
    -146.226130131271, -138.723605440997, 138.736376140396, 146.237519009027, 
    153.739441639357, 161.241995141072, 168.745010021227, 176.248305337399, 
    -176.248305337399, -168.745010021227, -161.241995141072, 
    -153.739441639357, -146.237519009027, -138.736376140396, 
    138.744789362256, 146.245184385179, 153.745894954228, 161.246868743795, 
    168.748039810838, 176.249332853807, -176.249332853807, -168.748039810838, 
    -161.246868743795, -153.745894954228, -146.245184385179, 
    -138.744789362256, 138.74895984555, 146.249033325085, 153.749171886272, 
    161.249365807297, 168.749601879962, 176.249864305626, -176.249864305626, 
    -168.749601879962, -161.249365807297, -153.749171886272, 
    -146.249033325085, -138.74895984555, 138.74895984555, 146.249033325085, 
    153.749171886272, 161.249365807297, 168.749601879962, 176.249864305626, 
    -176.249864305626, -168.749601879962, -161.249365807297, 
    -153.749171886272, -146.249033325085, -138.74895984555, 138.744789362256, 
    146.245184385179, 153.745894954228, 161.246868743795, 168.748039810838, 
    176.249332853807, -176.249332853807, -168.748039810838, 
    -161.246868743795, -153.745894954228, -146.245184385179, 
    -138.744789362256, 138.736376140396, 146.237519009027, 153.739441639357, 
    161.241995141072, 168.745010021227, 176.248305337399, -176.248305337399, 
    -168.745010021227, -161.241995141072, -153.739441639357, 
    -146.237519009027, -138.736376140396, 138.723605440997, 146.226130131271, 
    153.730028614144, 161.234988877032, 168.740697798093, 176.246850338243, 
    -176.246850338243, -168.740697798093, -161.234988877032, 
    -153.730028614144, -146.226130131271, -138.723605440997, 
    138.706389061519, 146.211228396465, 153.718017445191, 161.226220848091, 
    168.73537209375, 176.245065340346, -176.245065340346, -168.73537209375, 
    -161.226220848091, -153.718017445191, -146.211228396465, 
    -138.706389061519, 138.684791096902, 146.193228911696, 153.703950753707, 
    161.216189572235, 168.729373633571, 176.243070530866, -176.243070530866, 
    -168.729373633571, -161.216189572235, -153.703950753707, 
    -146.193228911696, -138.684791096902, -131.315208903098, 
    -123.806771088304, -116.296049246293, -108.783810427765, 
    -101.270626366429, -93.7569294691345, -86.2430705308655, 
    -78.7293736335712, -71.2161895722352, -63.7039507537071, 
    -56.193228911696, -48.6847910969017, -131.293610938481, 
    -123.788771603535, -116.281982554809, -108.773779151909, 
    -101.26462790625, -93.7549346596545, -86.2450653403455, 
    -78.7353720937503, -71.2262208480905, -63.7180174451908, 
    -56.2112283964646, -48.7063890615195, -131.276394559003, 
    -123.773869868729, -116.269971385856, -108.765011122968, 
    -101.259302201907, -93.7531496617566, -86.2468503382434, 
    -78.740697798093, -71.2349888770322, -63.7300286141441, -56.226130131271, 
    -48.7236054409966, -131.263623859604, -123.762480990973, 
    -116.260558360643, -108.758004858928, -101.254989978773, 
    -93.7516946626013, -86.2483053373987, -78.7450100212269, 
    -71.2419951410716, -63.7394416393566, -56.2375190090268, 
    -48.7363761403957, -131.255210637744, -123.754815614821, 
    -116.254105045772, -108.753131256205, -101.251960189162, 
    -93.7506671461934, -86.2493328538066, -78.7480398108377, 
    -71.2468687437952, -63.745894954228, -56.2451843851787, 
    -48.7447893622563, -131.25104015445, -123.750966674915, 
    -116.250828113728, -108.750634192703, -101.250398120038, 
    -93.7501356943742, -86.2498643056258, -78.7496018799618, 
    -71.2493658072972, -63.7491718862718, -56.2490333250849, 
    -48.7489598455498, -131.25104015445, -123.750966674915, 
    -116.250828113728, -108.750634192703, -101.250398120038, 
    -93.7501356943742, -86.2498643056258, -78.7496018799618, 
    -71.2493658072972, -63.7491718862718, -56.2490333250849, 
    -48.7489598455498, -131.255210637744, -123.754815614821, 
    -116.254105045772, -108.753131256205, -101.251960189162, 
    -93.7506671461934, -86.2493328538066, -78.7480398108377, 
    -71.2468687437952, -63.745894954228, -56.2451843851787, 
    -48.7447893622563, -131.263623859604, -123.762480990973, 
    -116.260558360643, -108.758004858928, -101.254989978773, 
    -93.7516946626013, -86.2483053373987, -78.7450100212268, 
    -71.2419951410716, -63.7394416393566, -56.2375190090268, 
    -48.7363761403957, -131.276394559003, -123.773869868729, 
    -116.269971385856, -108.765011122968, -101.259302201907, 
    -93.7531496617566, -86.2468503382434, -78.740697798093, 
    -71.2349888770322, -63.7300286141441, -56.226130131271, 
    -48.7236054409966, -131.293610938481, -123.788771603535, 
    -116.281982554809, -108.773779151909, -101.26462790625, 
    -93.7549346596545, -86.2450653403455, -78.7353720937503, 
    -71.2262208480905, -63.7180174451908, -56.2112283964646, 
    -48.7063890615195, -131.315208903098, -123.806771088304, 
    -116.296049246293, -108.783810427765, -101.270626366429, 
    -93.7569294691345, -86.2430705308655, -78.7293736335712, 
    -71.2161895722352, -63.7039507537071, -56.193228911696, 
    -48.6847910969017, -45, -52.6789833932524, -60.6230549375758, 
    -68.8117766657024, -77.1996324828867, -85.7180395939545, 
    -94.2819604060455, -102.800367517113, -111.188223334298, 
    -119.376945062424, -127.321016606748, -135, -37.3210166067476, -45, 
    -53.5572094377989, -63.0474748751433, -73.4040282512066, 
    -84.3904814032623, -95.6095185967377, -106.595971748793, 
    -116.952525124857, -126.442790562201, -135, -142.678983393252, 
    -29.3769450624242, -36.4427905622011, -45, -55.4480118954588, 
    -68.0198276783457, -82.4232160454614, -97.5767839545386, 
    -111.980172321654, -124.551988104541, -135, -143.557209437799, 
    -150.623054937576, -21.1882233342976, -26.9525251248567, 
    -34.5519881045412, -45, -59.6237942274726, -79.0670957284935, 
    -100.932904271507, -120.376205772527, -135, -145.448011895459, 
    -153.047474875143, -158.811776665702, -12.8003675171133, 
    -16.5959717487934, -21.9801723216543, -30.3762057725274, -45, 
    -71.7600509981516, -108.239949001848, -135, -149.623794227473, 
    -158.019827678346, -163.404028251207, -167.199632482887, 
    -4.28196040604547, -5.60951859673771, -7.57678395453862, 
    -10.9329042715065, -18.2399490018484, -45, -135, -161.760050998152, 
    -169.067095728493, -172.423216045461, -174.390481403262, 
    -175.718039593955, 4.28196040604546, 5.6095185967377, 7.57678395453862, 
    10.9329042715065, 18.2399490018484, 45, 135, 161.760050998152, 
    169.067095728493, 172.423216045461, 174.390481403262, 175.718039593955, 
    12.8003675171133, 16.5959717487934, 21.9801723216543, 30.3762057725274, 
    45, 71.7600509981516, 108.239949001848, 135, 149.623794227473, 
    158.019827678346, 163.404028251207, 167.199632482887, 21.1882233342975, 
    26.9525251248567, 34.5519881045412, 45, 59.6237942274726, 
    79.0670957284935, 100.932904271507, 120.376205772527, 135, 
    145.448011895459, 153.047474875143, 158.811776665702, 29.3769450624242, 
    36.4427905622011, 45, 55.4480118954588, 68.0198276783457, 
    82.4232160454614, 97.5767839545386, 111.980172321654, 124.551988104541, 
    135, 143.557209437799, 150.623054937576, 37.3210166067476, 45, 
    53.5572094377988, 63.0474748751433, 73.4040282512066, 84.3904814032623, 
    95.6095185967377, 106.595971748793, 116.952525124857, 126.442790562201, 
    135, 142.678983393252, 45, 52.6789833932524, 60.6230549375758, 
    68.8117766657024, 77.1996324828867, 85.7180395939545, 94.2819604060455, 
    102.800367517113, 111.188223334298, 119.376945062424, 127.321016606748, 
    135, 45, 52.6789833932524, 60.6230549375758, 68.8117766657024, 
    77.1996324828867, 85.7180395939545, 94.2819604060455, 102.800367517113, 
    111.188223334298, 119.376945062424, 127.321016606748, 135, 
    37.3210166067476, 45, 53.5572094377989, 63.0474748751433, 
    73.4040282512066, 84.3904814032623, 95.6095185967377, 106.595971748793, 
    116.952525124857, 126.442790562201, 135, 142.678983393252, 
    29.3769450624242, 36.4427905622011, 45, 55.4480118954588, 
    68.0198276783457, 82.4232160454614, 97.5767839545386, 111.980172321654, 
    124.551988104541, 135, 143.557209437799, 150.623054937576, 
    21.1882233342976, 26.9525251248567, 34.5519881045412, 45, 
    59.6237942274726, 79.0670957284935, 100.932904271507, 120.376205772527, 
    135, 145.448011895459, 153.047474875143, 158.811776665702, 
    12.8003675171133, 16.5959717487934, 21.9801723216543, 30.3762057725274, 
    45, 71.7600509981516, 108.239949001848, 135, 149.623794227473, 
    158.019827678346, 163.404028251207, 167.199632482887, 4.28196040604547, 
    5.60951859673771, 7.57678395453863, 10.9329042715065, 18.2399490018484, 
    45, 135, 161.760050998152, 169.067095728493, 172.423216045461, 
    174.390481403262, 175.718039593955, -4.28196040604547, -5.6095185967377, 
    -7.57678395453862, -10.9329042715065, -18.2399490018484, -45, -135, 
    -161.760050998152, -169.067095728493, -172.423216045461, 
    -174.390481403262, -175.718039593955, -12.8003675171133, 
    -16.5959717487934, -21.9801723216543, -30.3762057725274, -45, 
    -71.7600509981516, -108.239949001848, -135, -149.623794227473, 
    -158.019827678346, -163.404028251207, -167.199632482887, 
    -21.1882233342976, -26.9525251248567, -34.5519881045412, -45, 
    -59.6237942274726, -79.0670957284935, -100.932904271507, 
    -120.376205772527, -135, -145.448011895459, -153.047474875143, 
    -158.811776665702, -29.3769450624242, -36.4427905622011, -45, 
    -55.4480118954588, -68.0198276783457, -82.4232160454614, 
    -97.5767839545386, -111.980172321654, -124.551988104541, -135, 
    -143.557209437799, -150.623054937576, -37.3210166067476, -45, 
    -53.5572094377988, -63.0474748751433, -73.4040282512066, 
    -84.3904814032623, -95.6095185967377, -106.595971748793, 
    -116.952525124857, -126.442790562201, -135, -142.678983393252, -45, 
    -52.6789833932524, -60.6230549375758, -68.8117766657024, 
    -77.1996324828867, -85.7180395939545, -94.2819604060455, 
    -102.800367517113, -111.188223334298, -119.376945062424, 
    -127.321016606748, -135 ;

 dynamics_face_y = 33.432835056437, 36.1225579517621, 38.2011611172233, 
    39.7153031042524, 40.7028339742457, 41.1899453510804, 41.1899453510804, 
    40.7028339742457, 39.7153031042524, 38.2011611172233, 36.1225579517621, 
    33.432835056437, 26.7072135908547, 29.0798692007378, 30.9488663048686, 
    32.3308512179557, 33.2418639609319, 33.6941107346547, 33.6941107346547, 
    33.2418639609319, 32.3308512179557, 30.9488663048686, 29.0798692007378, 
    26.7072135908547, 20.3733724124488, 22.3180646012797, 23.8742427535654, 
    25.0396134449724, 25.8149813748506, 26.2020626588906, 26.2020626588906, 
    25.8149813748506, 25.0396134449724, 23.8742427535654, 22.3180646012797, 
    20.3733724124488, 14.3408794594474, 15.7797430199215, 16.9450166682866, 
    17.8263244005314, 18.417023334607, 18.7132512964975, 18.7132512964975, 
    18.417023334607, 17.8263244005314, 16.9450166682866, 15.7797430199215, 
    14.3408794594474, 8.52066086631705, 9.40290267273068, 10.1231569053278, 
    10.6715840982511, 11.0410464332339, 11.2269142890384, 11.2269142890384, 
    11.0410464332339, 10.6715840982511, 10.1231569053278, 9.40290267273068, 
    8.52066086631705, 2.82632454855766, 3.12345847186503, 3.36701515896158, 
    3.55310369075469, 3.67879389436188, 3.74212862554603, 3.74212862554603, 
    3.67879389436188, 3.55310369075469, 3.36701515896158, 3.12345847186503, 
    2.82632454855766, -2.82632454855766, -3.12345847186503, 
    -3.36701515896158, -3.55310369075468, -3.67879389436188, 
    -3.74212862554603, -3.74212862554603, -3.67879389436188, 
    -3.55310369075468, -3.36701515896158, -3.12345847186503, 
    -2.82632454855766, -8.52066086631705, -9.40290267273067, 
    -10.1231569053278, -10.6715840982511, -11.0410464332339, 
    -11.2269142890384, -11.2269142890384, -11.0410464332339, 
    -10.6715840982511, -10.1231569053278, -9.40290267273067, 
    -8.52066086631705, -14.3408794594474, -15.7797430199215, 
    -16.9450166682866, -17.8263244005314, -18.417023334607, 
    -18.7132512964974, -18.7132512964974, -18.417023334607, 
    -17.8263244005314, -16.9450166682866, -15.7797430199215, 
    -14.3408794594474, -20.3733724124488, -22.3180646012797, 
    -23.8742427535654, -25.0396134449724, -25.8149813748506, 
    -26.2020626588906, -26.2020626588906, -25.8149813748506, 
    -25.0396134449724, -23.8742427535654, -22.3180646012797, 
    -20.3733724124488, -26.7072135908547, -29.0798692007378, 
    -30.9488663048686, -32.3308512179557, -33.2418639609319, 
    -33.6941107346547, -33.6941107346547, -33.2418639609319, 
    -32.3308512179557, -30.9488663048686, -29.0798692007378, 
    -26.7072135908547, -33.432835056437, -36.1225579517621, 
    -38.2011611172233, -39.7153031042524, -40.7028339742457, 
    -41.1899453510804, -41.1899453510804, -40.7028339742457, 
    -39.7153031042524, -38.2011611172233, -36.1225579517621, 
    -33.432835056437, 33.432835056437, 36.1225579517621, 38.2011611172233, 
    39.7153031042524, 40.7028339742457, 41.1899453510804, 41.1899453510804, 
    40.7028339742457, 39.7153031042524, 38.2011611172233, 36.1225579517621, 
    33.432835056437, 26.7072135908547, 29.0798692007378, 30.9488663048686, 
    32.3308512179557, 33.2418639609319, 33.6941107346547, 33.6941107346547, 
    33.2418639609319, 32.3308512179557, 30.9488663048686, 29.0798692007378, 
    26.7072135908547, 20.3733724124488, 22.3180646012797, 23.8742427535654, 
    25.0396134449724, 25.8149813748506, 26.2020626588906, 26.2020626588906, 
    25.8149813748506, 25.0396134449724, 23.8742427535654, 22.3180646012797, 
    20.3733724124488, 14.3408794594474, 15.7797430199215, 16.9450166682866, 
    17.8263244005314, 18.417023334607, 18.7132512964975, 18.7132512964975, 
    18.417023334607, 17.8263244005314, 16.9450166682866, 15.7797430199215, 
    14.3408794594474, 8.52066086631705, 9.40290267273068, 10.1231569053278, 
    10.6715840982511, 11.0410464332339, 11.2269142890384, 11.2269142890384, 
    11.0410464332339, 10.6715840982511, 10.1231569053278, 9.40290267273068, 
    8.52066086631705, 2.82632454855766, 3.12345847186503, 3.36701515896158, 
    3.55310369075469, 3.67879389436188, 3.74212862554603, 3.74212862554603, 
    3.67879389436188, 3.55310369075469, 3.36701515896158, 3.12345847186503, 
    2.82632454855766, -2.82632454855766, -3.12345847186503, 
    -3.36701515896158, -3.55310369075468, -3.67879389436188, 
    -3.74212862554603, -3.74212862554603, -3.67879389436188, 
    -3.55310369075468, -3.36701515896158, -3.12345847186503, 
    -2.82632454855766, -8.52066086631705, -9.40290267273067, 
    -10.1231569053278, -10.6715840982511, -11.0410464332339, 
    -11.2269142890384, -11.2269142890384, -11.0410464332339, 
    -10.6715840982511, -10.1231569053278, -9.40290267273067, 
    -8.52066086631705, -14.3408794594474, -15.7797430199215, 
    -16.9450166682866, -17.8263244005314, -18.417023334607, 
    -18.7132512964974, -18.7132512964974, -18.417023334607, 
    -17.8263244005314, -16.9450166682866, -15.7797430199215, 
    -14.3408794594474, -20.3733724124488, -22.3180646012797, 
    -23.8742427535654, -25.0396134449724, -25.8149813748506, 
    -26.2020626588906, -26.2020626588906, -25.8149813748506, 
    -25.0396134449724, -23.8742427535654, -22.3180646012797, 
    -20.3733724124488, -26.7072135908547, -29.0798692007378, 
    -30.9488663048686, -32.3308512179557, -33.2418639609319, 
    -33.6941107346547, -33.6941107346547, -33.2418639609319, 
    -32.3308512179557, -30.9488663048686, -29.0798692007378, 
    -26.7072135908547, -33.432835056437, -36.1225579517621, 
    -38.2011611172233, -39.7153031042524, -40.7028339742457, 
    -41.1899453510804, -41.1899453510804, -40.7028339742457, 
    -39.7153031042524, -38.2011611172233, -36.1225579517621, 
    -33.432835056437, 33.432835056437, 36.1225579517621, 38.2011611172233, 
    39.7153031042524, 40.7028339742457, 41.1899453510804, 41.1899453510804, 
    40.7028339742457, 39.7153031042524, 38.2011611172233, 36.1225579517621, 
    33.432835056437, 26.7072135908547, 29.0798692007378, 30.9488663048686, 
    32.3308512179557, 33.2418639609319, 33.6941107346547, 33.6941107346547, 
    33.2418639609319, 32.3308512179557, 30.9488663048686, 29.0798692007378, 
    26.7072135908547, 20.3733724124488, 22.3180646012797, 23.8742427535654, 
    25.0396134449724, 25.8149813748506, 26.2020626588906, 26.2020626588906, 
    25.8149813748506, 25.0396134449724, 23.8742427535654, 22.3180646012797, 
    20.3733724124488, 14.3408794594474, 15.7797430199215, 16.9450166682866, 
    17.8263244005314, 18.417023334607, 18.7132512964975, 18.7132512964975, 
    18.417023334607, 17.8263244005314, 16.9450166682866, 15.7797430199215, 
    14.3408794594474, 8.52066086631705, 9.40290267273068, 10.1231569053278, 
    10.6715840982511, 11.0410464332339, 11.2269142890384, 11.2269142890384, 
    11.0410464332339, 10.6715840982511, 10.1231569053278, 9.40290267273068, 
    8.52066086631705, 2.82632454855766, 3.12345847186503, 3.36701515896158, 
    3.55310369075469, 3.67879389436188, 3.74212862554603, 3.74212862554603, 
    3.67879389436188, 3.55310369075469, 3.36701515896158, 3.12345847186503, 
    2.82632454855766, -2.82632454855766, -3.12345847186503, 
    -3.36701515896158, -3.55310369075468, -3.67879389436188, 
    -3.74212862554603, -3.74212862554603, -3.67879389436188, 
    -3.55310369075468, -3.36701515896158, -3.12345847186503, 
    -2.82632454855766, -8.52066086631705, -9.40290267273067, 
    -10.1231569053278, -10.6715840982511, -11.0410464332339, 
    -11.2269142890384, -11.2269142890384, -11.0410464332339, 
    -10.6715840982511, -10.1231569053278, -9.40290267273067, 
    -8.52066086631705, -14.3408794594474, -15.7797430199215, 
    -16.9450166682866, -17.8263244005314, -18.417023334607, 
    -18.7132512964974, -18.7132512964974, -18.417023334607, 
    -17.8263244005314, -16.9450166682866, -15.7797430199215, 
    -14.3408794594474, -20.3733724124488, -22.3180646012797, 
    -23.8742427535654, -25.0396134449724, -25.8149813748505, 
    -26.2020626588906, -26.2020626588906, -25.8149813748505, 
    -25.0396134449724, -23.8742427535654, -22.3180646012797, 
    -20.3733724124488, -26.7072135908547, -29.0798692007378, 
    -30.9488663048686, -32.3308512179557, -33.2418639609319, 
    -33.6941107346547, -33.6941107346547, -33.2418639609319, 
    -32.3308512179557, -30.9488663048686, -29.0798692007378, 
    -26.7072135908547, -33.432835056437, -36.1225579517621, 
    -38.2011611172233, -39.7153031042524, -40.7028339742457, 
    -41.1899453510804, -41.1899453510804, -40.7028339742457, 
    -39.7153031042524, -38.2011611172233, -36.1225579517621, 
    -33.432835056437, 33.432835056437, 36.1225579517621, 38.2011611172233, 
    39.7153031042524, 40.7028339742457, 41.1899453510804, 41.1899453510804, 
    40.7028339742457, 39.7153031042524, 38.2011611172233, 36.1225579517621, 
    33.432835056437, 26.7072135908547, 29.0798692007378, 30.9488663048686, 
    32.3308512179557, 33.2418639609319, 33.6941107346547, 33.6941107346547, 
    33.2418639609319, 32.3308512179557, 30.9488663048686, 29.0798692007378, 
    26.7072135908547, 20.3733724124488, 22.3180646012797, 23.8742427535654, 
    25.0396134449724, 25.8149813748506, 26.2020626588906, 26.2020626588906, 
    25.8149813748506, 25.0396134449724, 23.8742427535654, 22.3180646012797, 
    20.3733724124488, 14.3408794594474, 15.7797430199215, 16.9450166682866, 
    17.8263244005314, 18.417023334607, 18.7132512964975, 18.7132512964975, 
    18.417023334607, 17.8263244005314, 16.9450166682866, 15.7797430199215, 
    14.3408794594474, 8.52066086631705, 9.40290267273068, 10.1231569053278, 
    10.6715840982511, 11.0410464332339, 11.2269142890384, 11.2269142890384, 
    11.0410464332339, 10.6715840982511, 10.1231569053278, 9.40290267273068, 
    8.52066086631705, 2.82632454855766, 3.12345847186503, 3.36701515896158, 
    3.55310369075469, 3.67879389436188, 3.74212862554603, 3.74212862554603, 
    3.67879389436188, 3.55310369075469, 3.36701515896158, 3.12345847186503, 
    2.82632454855766, -2.82632454855766, -3.12345847186503, 
    -3.36701515896158, -3.55310369075468, -3.67879389436188, 
    -3.74212862554603, -3.74212862554603, -3.67879389436188, 
    -3.55310369075468, -3.36701515896158, -3.12345847186503, 
    -2.82632454855766, -8.52066086631705, -9.40290267273067, 
    -10.1231569053278, -10.6715840982511, -11.0410464332339, 
    -11.2269142890384, -11.2269142890384, -11.0410464332339, 
    -10.6715840982511, -10.1231569053278, -9.40290267273067, 
    -8.52066086631705, -14.3408794594474, -15.7797430199215, 
    -16.9450166682866, -17.8263244005314, -18.417023334607, 
    -18.7132512964974, -18.7132512964974, -18.417023334607, 
    -17.8263244005314, -16.9450166682866, -15.7797430199215, 
    -14.3408794594474, -20.3733724124488, -22.3180646012797, 
    -23.8742427535654, -25.0396134449724, -25.8149813748505, 
    -26.2020626588906, -26.2020626588906, -25.8149813748505, 
    -25.0396134449724, -23.8742427535654, -22.3180646012797, 
    -20.3733724124488, -26.7072135908547, -29.0798692007378, 
    -30.9488663048686, -32.3308512179557, -33.2418639609319, 
    -33.6941107346547, -33.6941107346547, -33.2418639609319, 
    -32.3308512179557, -30.9488663048686, -29.0798692007378, 
    -26.7072135908547, -33.432835056437, -36.1225579517621, 
    -38.2011611172233, -39.7153031042524, -40.7028339742457, 
    -41.1899453510804, -41.1899453510804, -40.7028339742457, 
    -39.7153031042524, -38.2011611172233, -36.1225579517621, 
    -33.432835056437, 38.8150077347025, 42.1582896974909, 44.7910057014103, 
    46.7407217209629, 48.028885464146, 48.6695532368043, 48.6695532368043, 
    48.028885464146, 46.7407217209629, 44.7910057014103, 42.1582896974909, 
    38.8150077347025, 42.1582896974908, 46.5794639642221, 50.2614918513234, 
    53.1318721567636, 55.1100100086019, 56.1218639580552, 56.1218639580552, 
    55.1100100086019, 53.1318721567636, 50.2614918513234, 46.5794639642222, 
    42.1582896974909, 44.7910057014103, 50.2614918513234, 55.083961998064, 
    59.0768040127068, 61.9916577943195, 63.5493286289719, 63.5493286289719, 
    61.9916577943195, 59.0768040127068, 55.083961998064, 50.2614918513234, 
    44.7910057014103, 46.7407217209629, 53.1318721567636, 59.0768040127068, 
    64.3459021628081, 68.5184407025596, 70.9275913731519, 70.9275913731519, 
    68.5184407025597, 64.3459021628081, 59.0768040127068, 53.1318721567636, 
    46.7407217209629, 48.028885464146, 55.1100100086019, 61.9916577943195, 
    68.5184407025597, 74.2857944271342, 78.1707754306064, 78.1707754306064, 
    74.2857944271342, 68.5184407025597, 61.9916577943196, 55.1100100086019, 
    48.028885464146, 48.6695532368043, 56.1218639580552, 63.5493286289719, 
    70.9275913731519, 78.1707754306064, 84.7040547607168, 84.7040547607168, 
    78.1707754306064, 70.9275913731519, 63.5493286289719, 56.1218639580552, 
    48.6695532368043, 48.6695532368043, 56.1218639580552, 63.5493286289719, 
    70.9275913731519, 78.1707754306064, 84.7040547607168, 84.7040547607168, 
    78.1707754306064, 70.9275913731519, 63.5493286289719, 56.1218639580552, 
    48.6695532368043, 48.028885464146, 55.1100100086019, 61.9916577943195, 
    68.5184407025597, 74.2857944271342, 78.1707754306064, 78.1707754306064, 
    74.2857944271342, 68.5184407025597, 61.9916577943196, 55.1100100086019, 
    48.028885464146, 46.7407217209629, 53.1318721567636, 59.0768040127068, 
    64.3459021628081, 68.5184407025597, 70.9275913731519, 70.9275913731519, 
    68.5184407025597, 64.3459021628081, 59.0768040127068, 53.1318721567636, 
    46.7407217209629, 44.7910057014103, 50.2614918513234, 55.083961998064, 
    59.0768040127068, 61.9916577943196, 63.5493286289719, 63.5493286289719, 
    61.9916577943196, 59.0768040127068, 55.083961998064, 50.2614918513234, 
    44.7910057014103, 42.1582896974909, 46.5794639642222, 50.2614918513234, 
    53.1318721567636, 55.1100100086019, 56.1218639580552, 56.1218639580552, 
    55.1100100086019, 53.1318721567636, 50.2614918513234, 46.5794639642222, 
    42.1582896974909, 38.8150077347025, 42.1582896974908, 44.7910057014103, 
    46.7407217209629, 48.028885464146, 48.6695532368043, 48.6695532368043, 
    48.028885464146, 46.7407217209629, 44.7910057014103, 42.1582896974909, 
    38.8150077347025, -38.8150077347025, -42.1582896974909, 
    -44.7910057014103, -46.7407217209629, -48.028885464146, 
    -48.6695532368043, -48.6695532368043, -48.028885464146, 
    -46.7407217209629, -44.7910057014103, -42.1582896974909, 
    -38.8150077347025, -42.1582896974909, -46.5794639642221, 
    -50.2614918513234, -53.1318721567636, -55.1100100086019, 
    -56.1218639580552, -56.1218639580552, -55.1100100086019, 
    -53.1318721567636, -50.2614918513234, -46.5794639642222, 
    -42.1582896974909, -44.7910057014103, -50.2614918513234, 
    -55.083961998064, -59.0768040127068, -61.9916577943195, 
    -63.5493286289719, -63.5493286289719, -61.9916577943195, 
    -59.0768040127068, -55.083961998064, -50.2614918513234, 
    -44.7910057014103, -46.7407217209629, -53.1318721567636, 
    -59.0768040127068, -64.3459021628081, -68.5184407025596, 
    -70.9275913731519, -70.9275913731519, -68.5184407025597, 
    -64.3459021628081, -59.0768040127068, -53.1318721567636, 
    -46.7407217209629, -48.028885464146, -55.1100100086019, 
    -61.9916577943195, -68.5184407025596, -74.2857944271342, 
    -78.1707754306064, -78.1707754306064, -74.2857944271342, 
    -68.5184407025597, -61.9916577943196, -55.1100100086019, 
    -48.028885464146, -48.6695532368043, -56.1218639580552, 
    -63.5493286289719, -70.9275913731519, -78.1707754306064, 
    -84.7040547607168, -84.7040547607168, -78.1707754306064, 
    -70.9275913731519, -63.5493286289719, -56.1218639580552, 
    -48.6695532368043, -48.6695532368043, -56.1218639580552, 
    -63.5493286289719, -70.9275913731519, -78.1707754306064, 
    -84.7040547607168, -84.7040547607168, -78.1707754306064, 
    -70.9275913731519, -63.5493286289719, -56.1218639580552, 
    -48.6695532368043, -48.028885464146, -55.1100100086019, 
    -61.9916577943195, -68.5184407025597, -74.2857944271342, 
    -78.1707754306064, -78.1707754306064, -74.2857944271342, 
    -68.5184407025597, -61.9916577943196, -55.1100100086019, 
    -48.028885464146, -46.7407217209629, -53.1318721567636, 
    -59.0768040127068, -64.3459021628081, -68.5184407025597, 
    -70.9275913731519, -70.9275913731519, -68.5184407025597, 
    -64.3459021628081, -59.0768040127068, -53.1318721567636, 
    -46.7407217209629, -44.7910057014103, -50.2614918513234, 
    -55.083961998064, -59.0768040127068, -61.9916577943196, 
    -63.5493286289719, -63.5493286289719, -61.9916577943196, 
    -59.0768040127068, -55.083961998064, -50.2614918513234, 
    -44.7910057014103, -42.1582896974909, -46.5794639642222, 
    -50.2614918513234, -53.1318721567636, -55.1100100086019, 
    -56.1218639580552, -56.1218639580552, -55.1100100086019, 
    -53.1318721567636, -50.2614918513234, -46.5794639642222, 
    -42.1582896974909, -38.8150077347025, -42.1582896974909, 
    -44.7910057014103, -46.7407217209629, -48.028885464146, 
    -48.6695532368043, -48.6695532368043, -48.028885464146, 
    -46.7407217209629, -44.7910057014103, -42.1582896974909, -38.8150077347025 ;
}
