netcdf split_file_2022121316-2022121320 {
dimensions:
	axis_nbounds = 2 ;
	lon = 1 ;
	lat = 1 ;
	nvertex = 2 ;
	levels = 39 ;
	time_counter = UNLIMITED ; // (5 currently)
variables:
	float lat(lat) ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:bounds = "bounds_lat" ;
	float lon(lon) ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:bounds = "bounds_lon" ;
	float bounds_lon(lat, lon, nvertex) ;
	float bounds_lat(lat, lon, nvertex) ;
	float levels(levels) ;
		levels:name = "levels" ;
		levels:units = "1" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 2022-12-13 01:00:00" ;
		time_instant:time_origin = "2022-12-13 01:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double time_counter(time_counter) ;
		time_counter:axis = "T" ;
		time_counter:standard_name = "time" ;
		time_counter:long_name = "Time axis" ;
		time_counter:calendar = "gregorian" ;
		time_counter:units = "seconds since 2022-12-13 01:00:00" ;
		time_counter:time_origin = "2022-12-13 01:00:00" ;
		time_counter:bounds = "time_counter_bounds" ;
	double time_counter_bounds(time_counter, axis_nbounds) ;
	float pressure(time_counter, levels, lat, lon) ;
		pressure:standard_name = "air_pressure" ;
		pressure:long_name = "Air Pressure" ;
		pressure:units = "Pa" ;
		pressure:online_operation = "instant" ;
		pressure:interval_operation = "1 h" ;
		pressure:interval_write = "1 h" ;
		pressure:cell_methods = "time: point" ;
		pressure:coordinates = "time_instant" ;
	float temperature(time_counter, levels, lat, lon) ;
		temperature:standard_name = "air_temperature" ;
		temperature:long_name = "Air Temperature" ;
		temperature:units = "K" ;
		temperature:online_operation = "instant" ;
		temperature:interval_operation = "1 h" ;
		temperature:interval_write = "1 h" ;
		temperature:cell_methods = "time: point" ;
		temperature:coordinates = "time_instant" ;

// global attributes:
		:name = "split_file" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "CF-1.6" ;
		:timeStamp = "2024-Jul-09 14:49:49 GMT" ;
		:uuid = "e4f7c26f-614c-43e1-8cea-4446ab4c92f8" ;
data:

 lat = 51.5 ;

 lon = -4.5 ;

 bounds_lon =
  -6, -3 ;

 bounds_lat =
  50, 53 ;

 levels = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 171, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39 ;

 time_instant = 57600, 61200, 64800, 68400, 72000 ;

 time_instant_bounds =
  57600, 57600,
  61200, 61200,
  64800, 64800,
  68400, 68400,
  72000, 72000 ;

 time_counter = 57600, 61200, 64800, 68400, 72000 ;

 time_counter_bounds =
  57600, 57600,
  61200, 61200,
  64800, 64800,
  68400, 68400,
  72000, 72000 ;

 pressure =
  1.609997e+07,
  1.609994e+07,
  1.609988e+07,
  1.609978e+07,
  1.609964e+07,
  1.609945e+07,
  1.609923e+07,
  1.609896e+07,
  1.609865e+07,
  1.60983e+07,
  1.609791e+07,
  1.609747e+07,
  1.609699e+07,
  1.609647e+07,
  1.60959e+07,
  1.609528e+07,
  1.609462e+07,
  1.60939e+07,
  1.609312e+07,
  1.609229e+07,
  1.609139e+07,
  1.609043e+07,
  1.60894e+07,
  1.608832e+07,
  1.608721e+07,
  1.608611e+07,
  1.6085e+07,
  1.608388e+07,
  1.608272e+07,
  1.608152e+07,
  1.608024e+07,
  1.607888e+07,
  1.607743e+07,
  1.607584e+07,
  1.607413e+07,
  1.607208e+07,
  1.606994e+07,
  1.606567e+07,
  1.606343e+07,
  1.709997e+07,
  1.709994e+07,
  1.709988e+07,
  1.709978e+07,
  1.709964e+07,
  1.709945e+07,
  1.709923e+07,
  1.709896e+07,
  1.709865e+07,
  1.70983e+07,
  1.709791e+07,
  1.709747e+07,
  1.709699e+07,
  1.709647e+07,
  1.70959e+07,
  1.709528e+07,
  1.709462e+07,
  1.70939e+07,
  1.709312e+07,
  1.709229e+07,
  1.709139e+07,
  1.709043e+07,
  1.70894e+07,
  1.708832e+07,
  1.708721e+07,
  1.708611e+07,
  1.7085e+07,
  1.708388e+07,
  1.708272e+07,
  1.708152e+07,
  1.708024e+07,
  1.707888e+07,
  1.707743e+07,
  1.707584e+07,
  1.707413e+07,
  1.707208e+07,
  1.706995e+07,
  1.706567e+07,
  1.706343e+07,
  1.809997e+07,
  1.809994e+07,
  1.809988e+07,
  1.809978e+07,
  1.809964e+07,
  1.809945e+07,
  1.809923e+07,
  1.809896e+07,
  1.809865e+07,
  1.80983e+07,
  1.809791e+07,
  1.809747e+07,
  1.809699e+07,
  1.809647e+07,
  1.80959e+07,
  1.809528e+07,
  1.809462e+07,
  1.80939e+07,
  1.809312e+07,
  1.809229e+07,
  1.809139e+07,
  1.809043e+07,
  1.80894e+07,
  1.808832e+07,
  1.808721e+07,
  1.808611e+07,
  1.8085e+07,
  1.808388e+07,
  1.808272e+07,
  1.808152e+07,
  1.808024e+07,
  1.807888e+07,
  1.807743e+07,
  1.807584e+07,
  1.807413e+07,
  1.807208e+07,
  1.806995e+07,
  1.806567e+07,
  1.806343e+07,
  1.909997e+07,
  1.909994e+07,
  1.909988e+07,
  1.909978e+07,
  1.909964e+07,
  1.909945e+07,
  1.909923e+07,
  1.909896e+07,
  1.909865e+07,
  1.90983e+07,
  1.909791e+07,
  1.909747e+07,
  1.909699e+07,
  1.909647e+07,
  1.90959e+07,
  1.909528e+07,
  1.909462e+07,
  1.90939e+07,
  1.909312e+07,
  1.909229e+07,
  1.909139e+07,
  1.909043e+07,
  1.90894e+07,
  1.908832e+07,
  1.908721e+07,
  1.908611e+07,
  1.9085e+07,
  1.908388e+07,
  1.908272e+07,
  1.908152e+07,
  1.908024e+07,
  1.907888e+07,
  1.907743e+07,
  1.907584e+07,
  1.907413e+07,
  1.907208e+07,
  1.906995e+07,
  1.906567e+07,
  1.906343e+07,
  2.009997e+07,
  2.009994e+07,
  2.009988e+07,
  2.009978e+07,
  2.009964e+07,
  2.009945e+07,
  2.009923e+07,
  2.009896e+07,
  2.009865e+07,
  2.00983e+07,
  2.009791e+07,
  2.009747e+07,
  2.009699e+07,
  2.009647e+07,
  2.00959e+07,
  2.009528e+07,
  2.009462e+07,
  2.00939e+07,
  2.009312e+07,
  2.009229e+07,
  2.009139e+07,
  2.009043e+07,
  2.00894e+07,
  2.008832e+07,
  2.008721e+07,
  2.008611e+07,
  2.0085e+07,
  2.008388e+07,
  2.008272e+07,
  2.008152e+07,
  2.008024e+07,
  2.007888e+07,
  2.007743e+07,
  2.007584e+07,
  2.007413e+07,
  2.007208e+07,
  2.006995e+07,
  2.006567e+07,
  2.006343e+07 ;

 temperature =
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600027e+07,
  1.600026e+07,
  1.600026e+07,
  1.600026e+07,
  1.600026e+07,
  1.600026e+07,
  1.600025e+07,
  1.600025e+07,
  1.600024e+07,
  1.600024e+07,
  1.600023e+07,
  1.600023e+07,
  1.600022e+07,
  1.600021e+07,
  1.600021e+07,
  1.600021e+07,
  1.600021e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600022e+07,
  1.600023e+07,
  1.600022e+07,
  1.600027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700027e+07,
  1.700026e+07,
  1.700026e+07,
  1.700026e+07,
  1.700026e+07,
  1.700025e+07,
  1.700025e+07,
  1.700024e+07,
  1.700024e+07,
  1.700023e+07,
  1.700023e+07,
  1.700022e+07,
  1.700021e+07,
  1.700021e+07,
  1.700021e+07,
  1.700021e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700022e+07,
  1.700023e+07,
  1.700022e+07,
  1.700027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800027e+07,
  1.800026e+07,
  1.800026e+07,
  1.800026e+07,
  1.800026e+07,
  1.800025e+07,
  1.800025e+07,
  1.800024e+07,
  1.800024e+07,
  1.800023e+07,
  1.800023e+07,
  1.800022e+07,
  1.800021e+07,
  1.800021e+07,
  1.800021e+07,
  1.800021e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800022e+07,
  1.800023e+07,
  1.800022e+07,
  1.800027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900027e+07,
  1.900026e+07,
  1.900026e+07,
  1.900026e+07,
  1.900026e+07,
  1.900025e+07,
  1.900025e+07,
  1.900024e+07,
  1.900024e+07,
  1.900023e+07,
  1.900023e+07,
  1.900022e+07,
  1.900021e+07,
  1.900021e+07,
  1.900021e+07,
  1.900021e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900022e+07,
  1.900023e+07,
  1.900022e+07,
  1.900027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000027e+07,
  2.000026e+07,
  2.000026e+07,
  2.000026e+07,
  2.000026e+07,
  2.000025e+07,
  2.000025e+07,
  2.000024e+07,
  2.000024e+07,
  2.000023e+07,
  2.000023e+07,
  2.000022e+07,
  2.000021e+07,
  2.000021e+07,
  2.000021e+07,
  2.000021e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000022e+07,
  2.000023e+07,
  2.000022e+07,
  2.000027e+07 ;
}
