netcdf domain_input {
dimensions:
        x = 5 ;
        y = 5 ;
variables:
        float x(x) ;
                x:long_name = "x coordinate" ;
                x:units = "1";
        float y(y) ;
                y:long_name = "y coordinate" ;
                y:units = "1";
        double field_A(y,x) ;
                field_A:long_name = "field A input data values" ;
                field_A:units = "1";

// global attributes:
                :title = "Field A input data" ;

data:

 x = 0, 2, 4, 6, 8 ;

 y = 0, 2, 4, 6, 8 ;


 field_A =  0,  4, 16, 36, 64,
                  4,  8, 20, 40, 68,
                 16, 20, 32, 52, 80,
                 36, 40, 52, 72, 100,
                 64, 68, 80, 100, 128 ;


}
